`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/27/2020 02:34:05 PM
// Design Name: 
// Module Name: asset
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module heart(
    (* synthesis, rom_block = "ROM_CELLXYZ01" *)
    input wire clk,
	input wire [3:0] x,
	input wire [3:0] y,
	output reg [11:0] rgb_reg
    );
    
    always @(posedge clk) begin
        case({y,x})
            8'b00000000: begin rgb_reg = 12'b000000000000; end
            8'b00000001: begin rgb_reg = 12'b000000000000; end
            8'b00000010: begin rgb_reg = 12'b000000000000; end
            8'b00000011: begin rgb_reg = 12'b000100010001; end
            8'b00000100: begin rgb_reg = 12'b000100010001; end
            8'b00000101: begin rgb_reg = 12'b000100010001; end
            8'b00000110: begin rgb_reg = 12'b000000000000; end
            8'b00000111: begin rgb_reg = 12'b000000000000; end
            8'b00001000: begin rgb_reg = 12'b000000000000; end
            8'b00001001: begin rgb_reg = 12'b000000000000; end
            8'b00001010: begin rgb_reg = 12'b000100010001; end
            8'b00001011: begin rgb_reg = 12'b000100010001; end
            8'b00001100: begin rgb_reg = 12'b000100010001; end
            8'b00001101: begin rgb_reg = 12'b000000000000; end
            8'b00001110: begin rgb_reg = 12'b000000000000; end
            8'b00001111: begin rgb_reg = 12'b000000000000; end
            8'b00010000: begin rgb_reg = 12'b000000000000; end
            8'b00010001: begin rgb_reg = 12'b000000000000; end
            8'b00010010: begin rgb_reg = 12'b000000000000; end
            8'b00010011: begin rgb_reg = 12'b010100010100; end
            8'b00010100: begin rgb_reg = 12'b011100100101; end
            8'b00010101: begin rgb_reg = 12'b011100100101; end
            8'b00010110: begin rgb_reg = 12'b000100010001; end
            8'b00010111: begin rgb_reg = 12'b000000000000; end
            8'b00011000: begin rgb_reg = 12'b000000000000; end
            8'b00011001: begin rgb_reg = 12'b000100010001; end
            8'b00011010: begin rgb_reg = 12'b011000100100; end
            8'b00011011: begin rgb_reg = 12'b011100100101; end
            8'b00011100: begin rgb_reg = 12'b011100100100; end
            8'b00011101: begin rgb_reg = 12'b000100010001; end
            8'b00011110: begin rgb_reg = 12'b000000000000; end
            8'b00011111: begin rgb_reg = 12'b000000000000; end
            8'b00100000: begin rgb_reg = 12'b000000000000; end
            8'b00100001: begin rgb_reg = 12'b000000010001; end
            8'b00100010: begin rgb_reg = 12'b011000100100; end
            8'b00100011: begin rgb_reg = 12'b110100000111; end
            8'b00100100: begin rgb_reg = 12'b111001001010; end
            8'b00100101: begin rgb_reg = 12'b111000011001; end
            8'b00100110: begin rgb_reg = 12'b100000010101; end
            8'b00100111: begin rgb_reg = 12'b001000010001; end
            8'b00101000: begin rgb_reg = 12'b000100010001; end
            8'b00101001: begin rgb_reg = 12'b011100100100; end
            8'b00101010: begin rgb_reg = 12'b111000000111; end
            8'b00101011: begin rgb_reg = 12'b111100001000; end
            8'b00101100: begin rgb_reg = 12'b111100000111; end
            8'b00101101: begin rgb_reg = 12'b011100100100; end
            8'b00101110: begin rgb_reg = 12'b000100010001; end
            8'b00101111: begin rgb_reg = 12'b000000000000; end
            8'b00110000: begin rgb_reg = 12'b000000010000; end
            8'b00110001: begin rgb_reg = 12'b011000010100; end
            8'b00110010: begin rgb_reg = 12'b111000001000; end
            8'b00110011: begin rgb_reg = 12'b111001001010; end
            8'b00110100: begin rgb_reg = 12'b111010001011; end
            8'b00110101: begin rgb_reg = 12'b111000101001; end
            8'b00110110: begin rgb_reg = 12'b111100001000; end
            8'b00110111: begin rgb_reg = 12'b100000010101; end
            8'b00111000: begin rgb_reg = 12'b011100100101; end
            8'b00111001: begin rgb_reg = 12'b111000001000; end
            8'b00111010: begin rgb_reg = 12'b111000000111; end
            8'b00111011: begin rgb_reg = 12'b111000001000; end
            8'b00111100: begin rgb_reg = 12'b111100001000; end
            8'b00111101: begin rgb_reg = 12'b111100000111; end
            8'b00111110: begin rgb_reg = 12'b011100100100; end
            8'b00111111: begin rgb_reg = 12'b000000010001; end
            8'b01000000: begin rgb_reg = 12'b001000110010; end
            8'b01000001: begin rgb_reg = 12'b110000000111; end
            8'b01000010: begin rgb_reg = 12'b111001011010; end
            8'b01000011: begin rgb_reg = 12'b111001111011; end
            8'b01000100: begin rgb_reg = 12'b111000011000; end
            8'b01000101: begin rgb_reg = 12'b111000000111; end
            8'b01000110: begin rgb_reg = 12'b111000000111; end
            8'b01000111: begin rgb_reg = 12'b111100001000; end
            8'b01001000: begin rgb_reg = 12'b111100001000; end
            8'b01001001: begin rgb_reg = 12'b111000000111; end
            8'b01001010: begin rgb_reg = 12'b111000000111; end
            8'b01001011: begin rgb_reg = 12'b111000000111; end
            8'b01001100: begin rgb_reg = 12'b111100001000; end
            8'b01001101: begin rgb_reg = 12'b111100000111; end
            8'b01001110: begin rgb_reg = 12'b111000000110; end
            8'b01001111: begin rgb_reg = 12'b001000110011; end
            8'b01010000: begin rgb_reg = 12'b001000110010; end
            8'b01010001: begin rgb_reg = 12'b110000000111; end
            8'b01010010: begin rgb_reg = 12'b111001111011; end
            8'b01010011: begin rgb_reg = 12'b111000011000; end
            8'b01010100: begin rgb_reg = 12'b111000000111; end
            8'b01010101: begin rgb_reg = 12'b111000000111; end
            8'b01010110: begin rgb_reg = 12'b111000000111; end
            8'b01010111: begin rgb_reg = 12'b111000000111; end
            8'b01011000: begin rgb_reg = 12'b111000000111; end
            8'b01011001: begin rgb_reg = 12'b111000000111; end
            8'b01011010: begin rgb_reg = 12'b111000000111; end
            8'b01011011: begin rgb_reg = 12'b111000000111; end
            8'b01011100: begin rgb_reg = 12'b111100001000; end
            8'b01011101: begin rgb_reg = 12'b111100000111; end
            8'b01011110: begin rgb_reg = 12'b111000000110; end
            8'b01011111: begin rgb_reg = 12'b001000110011; end
            8'b01100000: begin rgb_reg = 12'b001000110010; end
            8'b01100001: begin rgb_reg = 12'b110000000111; end
            8'b01100010: begin rgb_reg = 12'b111100001000; end
            8'b01100011: begin rgb_reg = 12'b111100001000; end
            8'b01100100: begin rgb_reg = 12'b111000000111; end
            8'b01100101: begin rgb_reg = 12'b111000000111; end
            8'b01100110: begin rgb_reg = 12'b111000000111; end
            8'b01100111: begin rgb_reg = 12'b111000000111; end
            8'b01101000: begin rgb_reg = 12'b111000000111; end
            8'b01101001: begin rgb_reg = 12'b111000000111; end
            8'b01101010: begin rgb_reg = 12'b111000000111; end
            8'b01101011: begin rgb_reg = 12'b111000000111; end
            8'b01101100: begin rgb_reg = 12'b111100001000; end
            8'b01101101: begin rgb_reg = 12'b111100000111; end
            8'b01101110: begin rgb_reg = 12'b111000000110; end
            8'b01101111: begin rgb_reg = 12'b001000110011; end
            8'b01110000: begin rgb_reg = 12'b000100010001; end
            8'b01110001: begin rgb_reg = 12'b100000010101; end
            8'b01110010: begin rgb_reg = 12'b111000000111; end
            8'b01110011: begin rgb_reg = 12'b111000000111; end
            8'b01110100: begin rgb_reg = 12'b111000000111; end
            8'b01110101: begin rgb_reg = 12'b111000000111; end
            8'b01110110: begin rgb_reg = 12'b111000000111; end
            8'b01110111: begin rgb_reg = 12'b111000000111; end
            8'b01111000: begin rgb_reg = 12'b111000000111; end
            8'b01111001: begin rgb_reg = 12'b111000000111; end
            8'b01111010: begin rgb_reg = 12'b111000000111; end
            8'b01111011: begin rgb_reg = 12'b111000001000; end
            8'b01111100: begin rgb_reg = 12'b111100000111; end
            8'b01111101: begin rgb_reg = 12'b111000000111; end
            8'b01111110: begin rgb_reg = 12'b100100010101; end
            8'b01111111: begin rgb_reg = 12'b000100010001; end
            8'b10000000: begin rgb_reg = 12'b000000000000; end
            8'b10000001: begin rgb_reg = 12'b001000100010; end
            8'b10000010: begin rgb_reg = 12'b110100000111; end
            8'b10000011: begin rgb_reg = 12'b111000000111; end
            8'b10000100: begin rgb_reg = 12'b111000000111; end
            8'b10000101: begin rgb_reg = 12'b111000000111; end
            8'b10000110: begin rgb_reg = 12'b111000000111; end
            8'b10000111: begin rgb_reg = 12'b111000000111; end
            8'b10001000: begin rgb_reg = 12'b111000000111; end
            8'b10001001: begin rgb_reg = 12'b111000000111; end
            8'b10001010: begin rgb_reg = 12'b111000000111; end
            8'b10001011: begin rgb_reg = 12'b111000000111; end
            8'b10001100: begin rgb_reg = 12'b111100000111; end
            8'b10001101: begin rgb_reg = 12'b111000000110; end
            8'b10001110: begin rgb_reg = 12'b001100110011; end
            8'b10001111: begin rgb_reg = 12'b000000000000; end
            8'b10010000: begin rgb_reg = 12'b000000000000; end
            8'b10010001: begin rgb_reg = 12'b000100010001; end
            8'b10010010: begin rgb_reg = 12'b100000010101; end
            8'b10010011: begin rgb_reg = 12'b110100000111; end
            8'b10010100: begin rgb_reg = 12'b111000000111; end
            8'b10010101: begin rgb_reg = 12'b111000000111; end
            8'b10010110: begin rgb_reg = 12'b111000000111; end
            8'b10010111: begin rgb_reg = 12'b111000000111; end
            8'b10011000: begin rgb_reg = 12'b111000000111; end
            8'b10011001: begin rgb_reg = 12'b111000000111; end
            8'b10011010: begin rgb_reg = 12'b111000000111; end
            8'b10011011: begin rgb_reg = 12'b111100000111; end
            8'b10011100: begin rgb_reg = 12'b111100000111; end
            8'b10011101: begin rgb_reg = 12'b100100010101; end
            8'b10011110: begin rgb_reg = 12'b000100010001; end
            8'b10011111: begin rgb_reg = 12'b000000000000; end
            8'b10100000: begin rgb_reg = 12'b000000000000; end
            8'b10100001: begin rgb_reg = 12'b000000000000; end
            8'b10100010: begin rgb_reg = 12'b000100010001; end
            8'b10100011: begin rgb_reg = 12'b011100010100; end
            8'b10100100: begin rgb_reg = 12'b111000000111; end
            8'b10100101: begin rgb_reg = 12'b111100000111; end
            8'b10100110: begin rgb_reg = 12'b111000000111; end
            8'b10100111: begin rgb_reg = 12'b111000000111; end
            8'b10101000: begin rgb_reg = 12'b111000000111; end
            8'b10101001: begin rgb_reg = 12'b111000000111; end
            8'b10101010: begin rgb_reg = 12'b111100000111; end
            8'b10101011: begin rgb_reg = 12'b111000000111; end
            8'b10101100: begin rgb_reg = 12'b101000010101; end
            8'b10101101: begin rgb_reg = 12'b000100010001; end
            8'b10101110: begin rgb_reg = 12'b000000000000; end
            8'b10101111: begin rgb_reg = 12'b000000000000; end
            8'b10110000: begin rgb_reg = 12'b000000000000; end
            8'b10110001: begin rgb_reg = 12'b000000000000; end
            8'b10110010: begin rgb_reg = 12'b000000000000; end
            8'b10110011: begin rgb_reg = 12'b000100010001; end
            8'b10110100: begin rgb_reg = 12'b100000010101; end
            8'b10110101: begin rgb_reg = 12'b110100000111; end
            8'b10110110: begin rgb_reg = 12'b111000001000; end
            8'b10110111: begin rgb_reg = 12'b111000000111; end
            8'b10111000: begin rgb_reg = 12'b111000000111; end
            8'b10111001: begin rgb_reg = 12'b111100000111; end
            8'b10111010: begin rgb_reg = 12'b111000000111; end
            8'b10111011: begin rgb_reg = 12'b100100010101; end
            8'b10111100: begin rgb_reg = 12'b001000010010; end
            8'b10111101: begin rgb_reg = 12'b000000000000; end
            8'b10111110: begin rgb_reg = 12'b000000000000; end
            8'b10111111: begin rgb_reg = 12'b000000000000; end
            8'b11000000: begin rgb_reg = 12'b000000000000; end
            8'b11000001: begin rgb_reg = 12'b000000000000; end
            8'b11000010: begin rgb_reg = 12'b000000000000; end
            8'b11000011: begin rgb_reg = 12'b000000000000; end
            8'b11000100: begin rgb_reg = 12'b000100010001; end
            8'b11000101: begin rgb_reg = 12'b011100010100; end
            8'b11000110: begin rgb_reg = 12'b111000000111; end
            8'b11000111: begin rgb_reg = 12'b111000001000; end
            8'b11001000: begin rgb_reg = 12'b111100000111; end
            8'b11001001: begin rgb_reg = 12'b111000000111; end
            8'b11001010: begin rgb_reg = 12'b100100010100; end
            8'b11001011: begin rgb_reg = 12'b000100010001; end
            8'b11001100: begin rgb_reg = 12'b000000000000; end
            8'b11001101: begin rgb_reg = 12'b000000000000; end
            8'b11001110: begin rgb_reg = 12'b000000000000; end
            8'b11001111: begin rgb_reg = 12'b000000000000; end
            8'b11010000: begin rgb_reg = 12'b000000000000; end
            8'b11010001: begin rgb_reg = 12'b000000000000; end
            8'b11010010: begin rgb_reg = 12'b000000000000; end
            8'b11010011: begin rgb_reg = 12'b000000000000; end
            8'b11010100: begin rgb_reg = 12'b000000000000; end
            8'b11010101: begin rgb_reg = 12'b000000010001; end
            8'b11010110: begin rgb_reg = 12'b100000010101; end
            8'b11010111: begin rgb_reg = 12'b111000000111; end
            8'b11011000: begin rgb_reg = 12'b111100000111; end
            8'b11011001: begin rgb_reg = 12'b100100010101; end
            8'b11011010: begin rgb_reg = 12'b001000100010; end
            8'b11011011: begin rgb_reg = 12'b000000000000; end
            8'b11011100: begin rgb_reg = 12'b000000000000; end
            8'b11011101: begin rgb_reg = 12'b000000000000; end
            8'b11011110: begin rgb_reg = 12'b000000000000; end
            8'b11011111: begin rgb_reg = 12'b000000000000; end
            8'b11100000: begin rgb_reg = 12'b000000000000; end
            8'b11100001: begin rgb_reg = 12'b000000000000; end
            8'b11100010: begin rgb_reg = 12'b000000000000; end
            8'b11100011: begin rgb_reg = 12'b000000000000; end
            8'b11100100: begin rgb_reg = 12'b000000000000; end
            8'b11100101: begin rgb_reg = 12'b000000000000; end
            8'b11100110: begin rgb_reg = 12'b000000010001; end
            8'b11100111: begin rgb_reg = 12'b100000010100; end
            8'b11101000: begin rgb_reg = 12'b100000010100; end
            8'b11101001: begin rgb_reg = 12'b000100010001; end
            8'b11101010: begin rgb_reg = 12'b000000000000; end
            8'b11101011: begin rgb_reg = 12'b000000000000; end
            8'b11101100: begin rgb_reg = 12'b000000000000; end
            8'b11101101: begin rgb_reg = 12'b000000000000; end
            8'b11101110: begin rgb_reg = 12'b000000000000; end
            8'b11101111: begin rgb_reg = 12'b000000000000; end
            8'b11110000: begin rgb_reg = 12'b000000000000; end
            8'b11110001: begin rgb_reg = 12'b000000000000; end
            8'b11110010: begin rgb_reg = 12'b000000000000; end
            8'b11110011: begin rgb_reg = 12'b000000000000; end
            8'b11110100: begin rgb_reg = 12'b000000000000; end
            8'b11110101: begin rgb_reg = 12'b000000000000; end
            8'b11110110: begin rgb_reg = 12'b000000000000; end
            8'b11110111: begin rgb_reg = 12'b000100010001; end
            8'b11111000: begin rgb_reg = 12'b000100010001; end
            8'b11111001: begin rgb_reg = 12'b000000000000; end
            8'b11111010: begin rgb_reg = 12'b000000000000; end
            8'b11111011: begin rgb_reg = 12'b000000000000; end
            8'b11111100: begin rgb_reg = 12'b000000000000; end
            8'b11111101: begin rgb_reg = 12'b000000000000; end
            8'b11111110: begin rgb_reg = 12'b000000000000; end
            8'b11111111: begin rgb_reg = 12'b000000000000; end
        endcase
    end  
endmodule

module menu(
    (* synthesis, rom_block = "ROM_CELLXYZ01" *)
    input wire clk,
	input wire [8:0] x,
	input wire [8:0] y,
	output reg [2:0] rgb_reg
    );
    
    always @(posedge clk) begin
        case({y,x})
            18'b000111000101101100: begin rgb_reg = 3'b001; end
            18'b000111000101101101: begin rgb_reg = 3'b011; end
            18'b000111000101101110: begin rgb_reg = 3'b011; end
            18'b000111000101101111: begin rgb_reg = 3'b011; end
            18'b000111000101110000: begin rgb_reg = 3'b011; end
            18'b000111000101110001: begin rgb_reg = 3'b011; end
            18'b000111000101110010: begin rgb_reg = 3'b011; end
            18'b000111000101110011: begin rgb_reg = 3'b011; end
            18'b000111000101110100: begin rgb_reg = 3'b011; end
            18'b000111001101101100: begin rgb_reg = 3'b001; end
            18'b000111001101101101: begin rgb_reg = 3'b001; end
            18'b000111001101101110: begin rgb_reg = 3'b001; end
            18'b000111001101101111: begin rgb_reg = 3'b001; end
            18'b000111001101110000: begin rgb_reg = 3'b001; end
            18'b000111001101110001: begin rgb_reg = 3'b001; end
            18'b000111001101110010: begin rgb_reg = 3'b001; end
            18'b000111001101110011: begin rgb_reg = 3'b001; end
            18'b000111001101110100: begin rgb_reg = 3'b001; end
            18'b000111010101101010: begin rgb_reg = 3'b001; end
            18'b000111010101101011: begin rgb_reg = 3'b011; end
            18'b000111010101110101: begin rgb_reg = 3'b011; end
            18'b000111010101110110: begin rgb_reg = 3'b001; end
            18'b000111011101101010: begin rgb_reg = 3'b001; end
            18'b000111011101101011: begin rgb_reg = 3'b011; end
            18'b000111011101110000: begin rgb_reg = 3'b001; end
            18'b000111011101110001: begin rgb_reg = 3'b001; end
            18'b000111011101110010: begin rgb_reg = 3'b001; end
            18'b000111011101110101: begin rgb_reg = 3'b011; end
            18'b000111011101110110: begin rgb_reg = 3'b001; end
            18'b000111100101101010: begin rgb_reg = 3'b001; end
            18'b000111100101101011: begin rgb_reg = 3'b011; end
            18'b000111100101110000: begin rgb_reg = 3'b011; end
            18'b000111100101110001: begin rgb_reg = 3'b011; end
            18'b000111100101110010: begin rgb_reg = 3'b011; end
            18'b000111100101110101: begin rgb_reg = 3'b011; end
            18'b000111100101110110: begin rgb_reg = 3'b001; end
            18'b000111101101101010: begin rgb_reg = 3'b001; end
            18'b000111101101101011: begin rgb_reg = 3'b011; end
            18'b000111101101101110: begin rgb_reg = 3'b001; end
            18'b000111101101101111: begin rgb_reg = 3'b001; end
            18'b000111101101110101: begin rgb_reg = 3'b011; end
            18'b000111101101110110: begin rgb_reg = 3'b001; end
            18'b000111110010011100: begin rgb_reg = 3'b001; end
            18'b000111110010011101: begin rgb_reg = 3'b011; end
            18'b000111110010011110: begin rgb_reg = 3'b011; end
            18'b000111110010011111: begin rgb_reg = 3'b011; end
            18'b000111110010101011: begin rgb_reg = 3'b001; end
            18'b000111110010101100: begin rgb_reg = 3'b011; end
            18'b000111110010101101: begin rgb_reg = 3'b011; end
            18'b000111110010101110: begin rgb_reg = 3'b011; end
            18'b000111110010110011: begin rgb_reg = 3'b011; end
            18'b000111110010110100: begin rgb_reg = 3'b011; end
            18'b000111110010110101: begin rgb_reg = 3'b011; end
            18'b000111110010110110: begin rgb_reg = 3'b011; end
            18'b000111110011000010: begin rgb_reg = 3'b011; end
            18'b000111110011000011: begin rgb_reg = 3'b011; end
            18'b000111110011000100: begin rgb_reg = 3'b011; end
            18'b000111110011000101: begin rgb_reg = 3'b011; end
            18'b000111110011001001: begin rgb_reg = 3'b001; end
            18'b000111110011001010: begin rgb_reg = 3'b011; end
            18'b000111110011001011: begin rgb_reg = 3'b011; end
            18'b000111110011001100: begin rgb_reg = 3'b011; end
            18'b000111110011001101: begin rgb_reg = 3'b011; end
            18'b000111110011001110: begin rgb_reg = 3'b011; end
            18'b000111110011001111: begin rgb_reg = 3'b011; end
            18'b000111110011010000: begin rgb_reg = 3'b011; end
            18'b000111110011010001: begin rgb_reg = 3'b011; end
            18'b000111110011010010: begin rgb_reg = 3'b011; end
            18'b000111110011010011: begin rgb_reg = 3'b011; end
            18'b000111110011010100: begin rgb_reg = 3'b011; end
            18'b000111110011010101: begin rgb_reg = 3'b011; end
            18'b000111110011010110: begin rgb_reg = 3'b011; end
            18'b000111110011010111: begin rgb_reg = 3'b011; end
            18'b000111110011011000: begin rgb_reg = 3'b001; end
            18'b000111110011100000: begin rgb_reg = 3'b011; end
            18'b000111110011100001: begin rgb_reg = 3'b011; end
            18'b000111110011100010: begin rgb_reg = 3'b011; end
            18'b000111110011100011: begin rgb_reg = 3'b011; end
            18'b000111110011100100: begin rgb_reg = 3'b011; end
            18'b000111110011100101: begin rgb_reg = 3'b011; end
            18'b000111110011100110: begin rgb_reg = 3'b011; end
            18'b000111110011100111: begin rgb_reg = 3'b011; end
            18'b000111110011101000: begin rgb_reg = 3'b011; end
            18'b000111110011101001: begin rgb_reg = 3'b011; end
            18'b000111110011101010: begin rgb_reg = 3'b011; end
            18'b000111110011101011: begin rgb_reg = 3'b011; end
            18'b000111110011101100: begin rgb_reg = 3'b011; end
            18'b000111110011101101: begin rgb_reg = 3'b011; end
            18'b000111110011101110: begin rgb_reg = 3'b011; end
            18'b000111110011101111: begin rgb_reg = 3'b011; end
            18'b000111110011110000: begin rgb_reg = 3'b011; end
            18'b000111110011110001: begin rgb_reg = 3'b011; end
            18'b000111110011110010: begin rgb_reg = 3'b011; end
            18'b000111110011110110: begin rgb_reg = 3'b001; end
            18'b000111110011110111: begin rgb_reg = 3'b011; end
            18'b000111110011111000: begin rgb_reg = 3'b011; end
            18'b000111110011111001: begin rgb_reg = 3'b011; end
            18'b000111110011111010: begin rgb_reg = 3'b011; end
            18'b000111110011111011: begin rgb_reg = 3'b011; end
            18'b000111110011111100: begin rgb_reg = 3'b011; end
            18'b000111110011111101: begin rgb_reg = 3'b011; end
            18'b000111110011111110: begin rgb_reg = 3'b011; end
            18'b000111110011111111: begin rgb_reg = 3'b011; end
            18'b000111110100000000: begin rgb_reg = 3'b011; end
            18'b000111110100000001: begin rgb_reg = 3'b011; end
            18'b000111110100000010: begin rgb_reg = 3'b011; end
            18'b000111110100000011: begin rgb_reg = 3'b011; end
            18'b000111110100000100: begin rgb_reg = 3'b011; end
            18'b000111110100000101: begin rgb_reg = 3'b001; end
            18'b000111110100001101: begin rgb_reg = 3'b011; end
            18'b000111110100001110: begin rgb_reg = 3'b011; end
            18'b000111110100001111: begin rgb_reg = 3'b011; end
            18'b000111110100010000: begin rgb_reg = 3'b011; end
            18'b000111110100011100: begin rgb_reg = 3'b011; end
            18'b000111110100011101: begin rgb_reg = 3'b011; end
            18'b000111110100011110: begin rgb_reg = 3'b011; end
            18'b000111110100011111: begin rgb_reg = 3'b011; end
            18'b000111110100100111: begin rgb_reg = 3'b011; end
            18'b000111110100101000: begin rgb_reg = 3'b011; end
            18'b000111110100101001: begin rgb_reg = 3'b011; end
            18'b000111110100101010: begin rgb_reg = 3'b011; end
            18'b000111110100101011: begin rgb_reg = 3'b011; end
            18'b000111110100101100: begin rgb_reg = 3'b011; end
            18'b000111110100101101: begin rgb_reg = 3'b011; end
            18'b000111110100101110: begin rgb_reg = 3'b011; end
            18'b000111110100101111: begin rgb_reg = 3'b011; end
            18'b000111110100110000: begin rgb_reg = 3'b011; end
            18'b000111110100110001: begin rgb_reg = 3'b011; end
            18'b000111110100110010: begin rgb_reg = 3'b001; end
            18'b000111110100111010: begin rgb_reg = 3'b011; end
            18'b000111110100111011: begin rgb_reg = 3'b011; end
            18'b000111110100111100: begin rgb_reg = 3'b011; end
            18'b000111110100111101: begin rgb_reg = 3'b011; end
            18'b000111110100111110: begin rgb_reg = 3'b011; end
            18'b000111110100111111: begin rgb_reg = 3'b011; end
            18'b000111110101000000: begin rgb_reg = 3'b011; end
            18'b000111110101000001: begin rgb_reg = 3'b011; end
            18'b000111110101000010: begin rgb_reg = 3'b011; end
            18'b000111110101000011: begin rgb_reg = 3'b011; end
            18'b000111110101000100: begin rgb_reg = 3'b011; end
            18'b000111110101000101: begin rgb_reg = 3'b011; end
            18'b000111110101000110: begin rgb_reg = 3'b011; end
            18'b000111110101000111: begin rgb_reg = 3'b011; end
            18'b000111110101001000: begin rgb_reg = 3'b011; end
            18'b000111110101010000: begin rgb_reg = 3'b001; end
            18'b000111110101010001: begin rgb_reg = 3'b011; end
            18'b000111110101010010: begin rgb_reg = 3'b011; end
            18'b000111110101010011: begin rgb_reg = 3'b011; end
            18'b000111110101010100: begin rgb_reg = 3'b011; end
            18'b000111110101010101: begin rgb_reg = 3'b011; end
            18'b000111110101010110: begin rgb_reg = 3'b011; end
            18'b000111110101010111: begin rgb_reg = 3'b011; end
            18'b000111110101011000: begin rgb_reg = 3'b011; end
            18'b000111110101011001: begin rgb_reg = 3'b011; end
            18'b000111110101011010: begin rgb_reg = 3'b011; end
            18'b000111110101011011: begin rgb_reg = 3'b011; end
            18'b000111110101011100: begin rgb_reg = 3'b011; end
            18'b000111110101011101: begin rgb_reg = 3'b011; end
            18'b000111110101011110: begin rgb_reg = 3'b011; end
            18'b000111110101011111: begin rgb_reg = 3'b011; end
            18'b000111110101100000: begin rgb_reg = 3'b011; end
            18'b000111110101100001: begin rgb_reg = 3'b011; end
            18'b000111110101100010: begin rgb_reg = 3'b011; end
            18'b000111110101101010: begin rgb_reg = 3'b001; end
            18'b000111110101101011: begin rgb_reg = 3'b011; end
            18'b000111110101101110: begin rgb_reg = 3'b011; end
            18'b000111110101101111: begin rgb_reg = 3'b001; end
            18'b000111110101110101: begin rgb_reg = 3'b011; end
            18'b000111110101110110: begin rgb_reg = 3'b001; end
            18'b000111111010011100: begin rgb_reg = 3'b001; end
            18'b000111111010011101: begin rgb_reg = 3'b011; end
            18'b000111111010011110: begin rgb_reg = 3'b011; end
            18'b000111111010011111: begin rgb_reg = 3'b011; end
            18'b000111111010101011: begin rgb_reg = 3'b001; end
            18'b000111111010101100: begin rgb_reg = 3'b011; end
            18'b000111111010101101: begin rgb_reg = 3'b011; end
            18'b000111111010101110: begin rgb_reg = 3'b011; end
            18'b000111111010110011: begin rgb_reg = 3'b011; end
            18'b000111111010110100: begin rgb_reg = 3'b011; end
            18'b000111111010110101: begin rgb_reg = 3'b011; end
            18'b000111111010110110: begin rgb_reg = 3'b011; end
            18'b000111111011000010: begin rgb_reg = 3'b011; end
            18'b000111111011000011: begin rgb_reg = 3'b011; end
            18'b000111111011000100: begin rgb_reg = 3'b011; end
            18'b000111111011000101: begin rgb_reg = 3'b011; end
            18'b000111111011001001: begin rgb_reg = 3'b001; end
            18'b000111111011001010: begin rgb_reg = 3'b011; end
            18'b000111111011001011: begin rgb_reg = 3'b011; end
            18'b000111111011001100: begin rgb_reg = 3'b011; end
            18'b000111111011001101: begin rgb_reg = 3'b011; end
            18'b000111111011001110: begin rgb_reg = 3'b011; end
            18'b000111111011001111: begin rgb_reg = 3'b011; end
            18'b000111111011010000: begin rgb_reg = 3'b011; end
            18'b000111111011010001: begin rgb_reg = 3'b011; end
            18'b000111111011010010: begin rgb_reg = 3'b011; end
            18'b000111111011010011: begin rgb_reg = 3'b011; end
            18'b000111111011010100: begin rgb_reg = 3'b011; end
            18'b000111111011010101: begin rgb_reg = 3'b011; end
            18'b000111111011010110: begin rgb_reg = 3'b011; end
            18'b000111111011010111: begin rgb_reg = 3'b011; end
            18'b000111111011011000: begin rgb_reg = 3'b001; end
            18'b000111111011100000: begin rgb_reg = 3'b011; end
            18'b000111111011100001: begin rgb_reg = 3'b011; end
            18'b000111111011100010: begin rgb_reg = 3'b011; end
            18'b000111111011100011: begin rgb_reg = 3'b011; end
            18'b000111111011100100: begin rgb_reg = 3'b011; end
            18'b000111111011100101: begin rgb_reg = 3'b011; end
            18'b000111111011100110: begin rgb_reg = 3'b011; end
            18'b000111111011100111: begin rgb_reg = 3'b011; end
            18'b000111111011101000: begin rgb_reg = 3'b011; end
            18'b000111111011101001: begin rgb_reg = 3'b011; end
            18'b000111111011101010: begin rgb_reg = 3'b011; end
            18'b000111111011101011: begin rgb_reg = 3'b011; end
            18'b000111111011101100: begin rgb_reg = 3'b011; end
            18'b000111111011101101: begin rgb_reg = 3'b011; end
            18'b000111111011101110: begin rgb_reg = 3'b011; end
            18'b000111111011101111: begin rgb_reg = 3'b011; end
            18'b000111111011110000: begin rgb_reg = 3'b011; end
            18'b000111111011110001: begin rgb_reg = 3'b011; end
            18'b000111111011110010: begin rgb_reg = 3'b011; end
            18'b000111111011110110: begin rgb_reg = 3'b001; end
            18'b000111111011110111: begin rgb_reg = 3'b011; end
            18'b000111111011111000: begin rgb_reg = 3'b011; end
            18'b000111111011111001: begin rgb_reg = 3'b011; end
            18'b000111111011111010: begin rgb_reg = 3'b011; end
            18'b000111111011111011: begin rgb_reg = 3'b011; end
            18'b000111111011111100: begin rgb_reg = 3'b011; end
            18'b000111111011111101: begin rgb_reg = 3'b011; end
            18'b000111111011111110: begin rgb_reg = 3'b011; end
            18'b000111111011111111: begin rgb_reg = 3'b011; end
            18'b000111111100000000: begin rgb_reg = 3'b011; end
            18'b000111111100000001: begin rgb_reg = 3'b011; end
            18'b000111111100000010: begin rgb_reg = 3'b011; end
            18'b000111111100000011: begin rgb_reg = 3'b011; end
            18'b000111111100000100: begin rgb_reg = 3'b011; end
            18'b000111111100000101: begin rgb_reg = 3'b001; end
            18'b000111111100001101: begin rgb_reg = 3'b011; end
            18'b000111111100001110: begin rgb_reg = 3'b011; end
            18'b000111111100001111: begin rgb_reg = 3'b011; end
            18'b000111111100010000: begin rgb_reg = 3'b011; end
            18'b000111111100011100: begin rgb_reg = 3'b011; end
            18'b000111111100011101: begin rgb_reg = 3'b011; end
            18'b000111111100011110: begin rgb_reg = 3'b011; end
            18'b000111111100011111: begin rgb_reg = 3'b011; end
            18'b000111111100100111: begin rgb_reg = 3'b011; end
            18'b000111111100101000: begin rgb_reg = 3'b011; end
            18'b000111111100101001: begin rgb_reg = 3'b011; end
            18'b000111111100101010: begin rgb_reg = 3'b011; end
            18'b000111111100101011: begin rgb_reg = 3'b011; end
            18'b000111111100101100: begin rgb_reg = 3'b011; end
            18'b000111111100101101: begin rgb_reg = 3'b011; end
            18'b000111111100101110: begin rgb_reg = 3'b011; end
            18'b000111111100101111: begin rgb_reg = 3'b011; end
            18'b000111111100110000: begin rgb_reg = 3'b011; end
            18'b000111111100110001: begin rgb_reg = 3'b011; end
            18'b000111111100110010: begin rgb_reg = 3'b001; end
            18'b000111111100111010: begin rgb_reg = 3'b011; end
            18'b000111111100111011: begin rgb_reg = 3'b011; end
            18'b000111111100111100: begin rgb_reg = 3'b011; end
            18'b000111111100111101: begin rgb_reg = 3'b011; end
            18'b000111111100111110: begin rgb_reg = 3'b011; end
            18'b000111111100111111: begin rgb_reg = 3'b011; end
            18'b000111111101000000: begin rgb_reg = 3'b011; end
            18'b000111111101000001: begin rgb_reg = 3'b011; end
            18'b000111111101000010: begin rgb_reg = 3'b011; end
            18'b000111111101000011: begin rgb_reg = 3'b011; end
            18'b000111111101000100: begin rgb_reg = 3'b011; end
            18'b000111111101000101: begin rgb_reg = 3'b011; end
            18'b000111111101000110: begin rgb_reg = 3'b011; end
            18'b000111111101000111: begin rgb_reg = 3'b011; end
            18'b000111111101001000: begin rgb_reg = 3'b011; end
            18'b000111111101010000: begin rgb_reg = 3'b001; end
            18'b000111111101010001: begin rgb_reg = 3'b011; end
            18'b000111111101010010: begin rgb_reg = 3'b011; end
            18'b000111111101010011: begin rgb_reg = 3'b011; end
            18'b000111111101010100: begin rgb_reg = 3'b011; end
            18'b000111111101010101: begin rgb_reg = 3'b011; end
            18'b000111111101010110: begin rgb_reg = 3'b011; end
            18'b000111111101010111: begin rgb_reg = 3'b011; end
            18'b000111111101011000: begin rgb_reg = 3'b011; end
            18'b000111111101011001: begin rgb_reg = 3'b011; end
            18'b000111111101011010: begin rgb_reg = 3'b011; end
            18'b000111111101011011: begin rgb_reg = 3'b011; end
            18'b000111111101011100: begin rgb_reg = 3'b011; end
            18'b000111111101011101: begin rgb_reg = 3'b011; end
            18'b000111111101011110: begin rgb_reg = 3'b011; end
            18'b000111111101011111: begin rgb_reg = 3'b011; end
            18'b000111111101100000: begin rgb_reg = 3'b011; end
            18'b000111111101100001: begin rgb_reg = 3'b011; end
            18'b000111111101100010: begin rgb_reg = 3'b011; end
            18'b000111111101101010: begin rgb_reg = 3'b001; end
            18'b000111111101101011: begin rgb_reg = 3'b011; end
            18'b000111111101110000: begin rgb_reg = 3'b011; end
            18'b000111111101110001: begin rgb_reg = 3'b011; end
            18'b000111111101110010: begin rgb_reg = 3'b011; end
            18'b000111111101110101: begin rgb_reg = 3'b011; end
            18'b000111111101110110: begin rgb_reg = 3'b001; end
            18'b001000000010011100: begin rgb_reg = 3'b001; end
            18'b001000000010011101: begin rgb_reg = 3'b011; end
            18'b001000000010011110: begin rgb_reg = 3'b011; end
            18'b001000000010011111: begin rgb_reg = 3'b011; end
            18'b001000000010101011: begin rgb_reg = 3'b001; end
            18'b001000000010101100: begin rgb_reg = 3'b011; end
            18'b001000000010101101: begin rgb_reg = 3'b011; end
            18'b001000000010101110: begin rgb_reg = 3'b011; end
            18'b001000000010110011: begin rgb_reg = 3'b011; end
            18'b001000000010110100: begin rgb_reg = 3'b011; end
            18'b001000000010110101: begin rgb_reg = 3'b011; end
            18'b001000000010110110: begin rgb_reg = 3'b011; end
            18'b001000000011000010: begin rgb_reg = 3'b011; end
            18'b001000000011000011: begin rgb_reg = 3'b011; end
            18'b001000000011000100: begin rgb_reg = 3'b011; end
            18'b001000000011000101: begin rgb_reg = 3'b011; end
            18'b001000000011001001: begin rgb_reg = 3'b001; end
            18'b001000000011001010: begin rgb_reg = 3'b011; end
            18'b001000000011001011: begin rgb_reg = 3'b011; end
            18'b001000000011001100: begin rgb_reg = 3'b011; end
            18'b001000000011001101: begin rgb_reg = 3'b011; end
            18'b001000000011001110: begin rgb_reg = 3'b011; end
            18'b001000000011001111: begin rgb_reg = 3'b011; end
            18'b001000000011010000: begin rgb_reg = 3'b011; end
            18'b001000000011010001: begin rgb_reg = 3'b011; end
            18'b001000000011010010: begin rgb_reg = 3'b011; end
            18'b001000000011010011: begin rgb_reg = 3'b011; end
            18'b001000000011010100: begin rgb_reg = 3'b011; end
            18'b001000000011010101: begin rgb_reg = 3'b011; end
            18'b001000000011010110: begin rgb_reg = 3'b011; end
            18'b001000000011010111: begin rgb_reg = 3'b011; end
            18'b001000000011011000: begin rgb_reg = 3'b001; end
            18'b001000000011100000: begin rgb_reg = 3'b011; end
            18'b001000000011100001: begin rgb_reg = 3'b011; end
            18'b001000000011100010: begin rgb_reg = 3'b011; end
            18'b001000000011100011: begin rgb_reg = 3'b011; end
            18'b001000000011100100: begin rgb_reg = 3'b011; end
            18'b001000000011100101: begin rgb_reg = 3'b011; end
            18'b001000000011100110: begin rgb_reg = 3'b011; end
            18'b001000000011100111: begin rgb_reg = 3'b011; end
            18'b001000000011101000: begin rgb_reg = 3'b011; end
            18'b001000000011101001: begin rgb_reg = 3'b011; end
            18'b001000000011101010: begin rgb_reg = 3'b011; end
            18'b001000000011101011: begin rgb_reg = 3'b011; end
            18'b001000000011101100: begin rgb_reg = 3'b011; end
            18'b001000000011101101: begin rgb_reg = 3'b011; end
            18'b001000000011101110: begin rgb_reg = 3'b011; end
            18'b001000000011101111: begin rgb_reg = 3'b011; end
            18'b001000000011110000: begin rgb_reg = 3'b011; end
            18'b001000000011110001: begin rgb_reg = 3'b011; end
            18'b001000000011110010: begin rgb_reg = 3'b011; end
            18'b001000000011110110: begin rgb_reg = 3'b001; end
            18'b001000000011110111: begin rgb_reg = 3'b011; end
            18'b001000000011111000: begin rgb_reg = 3'b011; end
            18'b001000000011111001: begin rgb_reg = 3'b011; end
            18'b001000000011111010: begin rgb_reg = 3'b011; end
            18'b001000000011111011: begin rgb_reg = 3'b011; end
            18'b001000000011111100: begin rgb_reg = 3'b011; end
            18'b001000000011111101: begin rgb_reg = 3'b011; end
            18'b001000000011111110: begin rgb_reg = 3'b011; end
            18'b001000000011111111: begin rgb_reg = 3'b011; end
            18'b001000000100000000: begin rgb_reg = 3'b011; end
            18'b001000000100000001: begin rgb_reg = 3'b011; end
            18'b001000000100000010: begin rgb_reg = 3'b011; end
            18'b001000000100000011: begin rgb_reg = 3'b011; end
            18'b001000000100000100: begin rgb_reg = 3'b011; end
            18'b001000000100000101: begin rgb_reg = 3'b001; end
            18'b001000000100001101: begin rgb_reg = 3'b011; end
            18'b001000000100001110: begin rgb_reg = 3'b011; end
            18'b001000000100001111: begin rgb_reg = 3'b011; end
            18'b001000000100010000: begin rgb_reg = 3'b011; end
            18'b001000000100011100: begin rgb_reg = 3'b011; end
            18'b001000000100011101: begin rgb_reg = 3'b011; end
            18'b001000000100011110: begin rgb_reg = 3'b011; end
            18'b001000000100011111: begin rgb_reg = 3'b011; end
            18'b001000000100100111: begin rgb_reg = 3'b011; end
            18'b001000000100101000: begin rgb_reg = 3'b011; end
            18'b001000000100101001: begin rgb_reg = 3'b011; end
            18'b001000000100101010: begin rgb_reg = 3'b011; end
            18'b001000000100101011: begin rgb_reg = 3'b011; end
            18'b001000000100101100: begin rgb_reg = 3'b011; end
            18'b001000000100101101: begin rgb_reg = 3'b011; end
            18'b001000000100101110: begin rgb_reg = 3'b011; end
            18'b001000000100101111: begin rgb_reg = 3'b011; end
            18'b001000000100110000: begin rgb_reg = 3'b011; end
            18'b001000000100110001: begin rgb_reg = 3'b011; end
            18'b001000000100110010: begin rgb_reg = 3'b001; end
            18'b001000000100111010: begin rgb_reg = 3'b011; end
            18'b001000000100111011: begin rgb_reg = 3'b011; end
            18'b001000000100111100: begin rgb_reg = 3'b011; end
            18'b001000000100111101: begin rgb_reg = 3'b011; end
            18'b001000000100111110: begin rgb_reg = 3'b011; end
            18'b001000000100111111: begin rgb_reg = 3'b011; end
            18'b001000000101000000: begin rgb_reg = 3'b011; end
            18'b001000000101000001: begin rgb_reg = 3'b011; end
            18'b001000000101000010: begin rgb_reg = 3'b011; end
            18'b001000000101000011: begin rgb_reg = 3'b011; end
            18'b001000000101000100: begin rgb_reg = 3'b011; end
            18'b001000000101000101: begin rgb_reg = 3'b011; end
            18'b001000000101000110: begin rgb_reg = 3'b011; end
            18'b001000000101000111: begin rgb_reg = 3'b011; end
            18'b001000000101001000: begin rgb_reg = 3'b011; end
            18'b001000000101010000: begin rgb_reg = 3'b001; end
            18'b001000000101010001: begin rgb_reg = 3'b011; end
            18'b001000000101010010: begin rgb_reg = 3'b011; end
            18'b001000000101010011: begin rgb_reg = 3'b011; end
            18'b001000000101010100: begin rgb_reg = 3'b011; end
            18'b001000000101010101: begin rgb_reg = 3'b011; end
            18'b001000000101010110: begin rgb_reg = 3'b011; end
            18'b001000000101010111: begin rgb_reg = 3'b011; end
            18'b001000000101011000: begin rgb_reg = 3'b011; end
            18'b001000000101011001: begin rgb_reg = 3'b011; end
            18'b001000000101011010: begin rgb_reg = 3'b011; end
            18'b001000000101011011: begin rgb_reg = 3'b011; end
            18'b001000000101011100: begin rgb_reg = 3'b011; end
            18'b001000000101011101: begin rgb_reg = 3'b011; end
            18'b001000000101011110: begin rgb_reg = 3'b011; end
            18'b001000000101011111: begin rgb_reg = 3'b011; end
            18'b001000000101100000: begin rgb_reg = 3'b011; end
            18'b001000000101100001: begin rgb_reg = 3'b011; end
            18'b001000000101100010: begin rgb_reg = 3'b011; end
            18'b001000000101101010: begin rgb_reg = 3'b001; end
            18'b001000000101101011: begin rgb_reg = 3'b011; end
            18'b001000000101110000: begin rgb_reg = 3'b001; end
            18'b001000000101110001: begin rgb_reg = 3'b001; end
            18'b001000000101110010: begin rgb_reg = 3'b001; end
            18'b001000000101110101: begin rgb_reg = 3'b011; end
            18'b001000000101110110: begin rgb_reg = 3'b001; end
            18'b001000001010011100: begin rgb_reg = 3'b001; end
            18'b001000001010011101: begin rgb_reg = 3'b011; end
            18'b001000001010011110: begin rgb_reg = 3'b011; end
            18'b001000001010011111: begin rgb_reg = 3'b011; end
            18'b001000001010101011: begin rgb_reg = 3'b001; end
            18'b001000001010101100: begin rgb_reg = 3'b011; end
            18'b001000001010101101: begin rgb_reg = 3'b011; end
            18'b001000001010101110: begin rgb_reg = 3'b011; end
            18'b001000001010110011: begin rgb_reg = 3'b011; end
            18'b001000001010110100: begin rgb_reg = 3'b011; end
            18'b001000001010110101: begin rgb_reg = 3'b011; end
            18'b001000001010110110: begin rgb_reg = 3'b011; end
            18'b001000001011000010: begin rgb_reg = 3'b011; end
            18'b001000001011000011: begin rgb_reg = 3'b011; end
            18'b001000001011000100: begin rgb_reg = 3'b011; end
            18'b001000001011000101: begin rgb_reg = 3'b011; end
            18'b001000001011001001: begin rgb_reg = 3'b001; end
            18'b001000001011001010: begin rgb_reg = 3'b011; end
            18'b001000001011001011: begin rgb_reg = 3'b011; end
            18'b001000001011001100: begin rgb_reg = 3'b011; end
            18'b001000001011001101: begin rgb_reg = 3'b011; end
            18'b001000001011001110: begin rgb_reg = 3'b011; end
            18'b001000001011001111: begin rgb_reg = 3'b011; end
            18'b001000001011010000: begin rgb_reg = 3'b011; end
            18'b001000001011010001: begin rgb_reg = 3'b011; end
            18'b001000001011010010: begin rgb_reg = 3'b011; end
            18'b001000001011010011: begin rgb_reg = 3'b011; end
            18'b001000001011010100: begin rgb_reg = 3'b011; end
            18'b001000001011010101: begin rgb_reg = 3'b011; end
            18'b001000001011010110: begin rgb_reg = 3'b011; end
            18'b001000001011010111: begin rgb_reg = 3'b011; end
            18'b001000001011011000: begin rgb_reg = 3'b001; end
            18'b001000001011100000: begin rgb_reg = 3'b011; end
            18'b001000001011100001: begin rgb_reg = 3'b011; end
            18'b001000001011100010: begin rgb_reg = 3'b011; end
            18'b001000001011100011: begin rgb_reg = 3'b011; end
            18'b001000001011100100: begin rgb_reg = 3'b011; end
            18'b001000001011100101: begin rgb_reg = 3'b011; end
            18'b001000001011100110: begin rgb_reg = 3'b011; end
            18'b001000001011100111: begin rgb_reg = 3'b011; end
            18'b001000001011101000: begin rgb_reg = 3'b011; end
            18'b001000001011101001: begin rgb_reg = 3'b011; end
            18'b001000001011101010: begin rgb_reg = 3'b011; end
            18'b001000001011101011: begin rgb_reg = 3'b011; end
            18'b001000001011101100: begin rgb_reg = 3'b011; end
            18'b001000001011101101: begin rgb_reg = 3'b011; end
            18'b001000001011101110: begin rgb_reg = 3'b011; end
            18'b001000001011101111: begin rgb_reg = 3'b011; end
            18'b001000001011110000: begin rgb_reg = 3'b011; end
            18'b001000001011110001: begin rgb_reg = 3'b011; end
            18'b001000001011110010: begin rgb_reg = 3'b001; end
            18'b001000001011110110: begin rgb_reg = 3'b001; end
            18'b001000001011110111: begin rgb_reg = 3'b011; end
            18'b001000001011111000: begin rgb_reg = 3'b011; end
            18'b001000001011111001: begin rgb_reg = 3'b011; end
            18'b001000001011111010: begin rgb_reg = 3'b011; end
            18'b001000001011111011: begin rgb_reg = 3'b011; end
            18'b001000001011111100: begin rgb_reg = 3'b011; end
            18'b001000001011111101: begin rgb_reg = 3'b011; end
            18'b001000001011111110: begin rgb_reg = 3'b011; end
            18'b001000001011111111: begin rgb_reg = 3'b011; end
            18'b001000001100000000: begin rgb_reg = 3'b011; end
            18'b001000001100000001: begin rgb_reg = 3'b011; end
            18'b001000001100000010: begin rgb_reg = 3'b011; end
            18'b001000001100000011: begin rgb_reg = 3'b011; end
            18'b001000001100000100: begin rgb_reg = 3'b011; end
            18'b001000001100000101: begin rgb_reg = 3'b001; end
            18'b001000001100001101: begin rgb_reg = 3'b011; end
            18'b001000001100001110: begin rgb_reg = 3'b011; end
            18'b001000001100001111: begin rgb_reg = 3'b011; end
            18'b001000001100010000: begin rgb_reg = 3'b011; end
            18'b001000001100011100: begin rgb_reg = 3'b011; end
            18'b001000001100011101: begin rgb_reg = 3'b011; end
            18'b001000001100011110: begin rgb_reg = 3'b011; end
            18'b001000001100011111: begin rgb_reg = 3'b011; end
            18'b001000001100100111: begin rgb_reg = 3'b001; end
            18'b001000001100101000: begin rgb_reg = 3'b011; end
            18'b001000001100101001: begin rgb_reg = 3'b011; end
            18'b001000001100101010: begin rgb_reg = 3'b011; end
            18'b001000001100101011: begin rgb_reg = 3'b011; end
            18'b001000001100101100: begin rgb_reg = 3'b011; end
            18'b001000001100101101: begin rgb_reg = 3'b011; end
            18'b001000001100101110: begin rgb_reg = 3'b011; end
            18'b001000001100101111: begin rgb_reg = 3'b011; end
            18'b001000001100110000: begin rgb_reg = 3'b011; end
            18'b001000001100110001: begin rgb_reg = 3'b011; end
            18'b001000001100110010: begin rgb_reg = 3'b001; end
            18'b001000001100111010: begin rgb_reg = 3'b011; end
            18'b001000001100111011: begin rgb_reg = 3'b011; end
            18'b001000001100111100: begin rgb_reg = 3'b011; end
            18'b001000001100111101: begin rgb_reg = 3'b011; end
            18'b001000001100111110: begin rgb_reg = 3'b011; end
            18'b001000001100111111: begin rgb_reg = 3'b011; end
            18'b001000001101000000: begin rgb_reg = 3'b011; end
            18'b001000001101000001: begin rgb_reg = 3'b011; end
            18'b001000001101000010: begin rgb_reg = 3'b011; end
            18'b001000001101000011: begin rgb_reg = 3'b011; end
            18'b001000001101000100: begin rgb_reg = 3'b011; end
            18'b001000001101000101: begin rgb_reg = 3'b011; end
            18'b001000001101000110: begin rgb_reg = 3'b011; end
            18'b001000001101000111: begin rgb_reg = 3'b011; end
            18'b001000001101001000: begin rgb_reg = 3'b011; end
            18'b001000001101010000: begin rgb_reg = 3'b001; end
            18'b001000001101010001: begin rgb_reg = 3'b011; end
            18'b001000001101010010: begin rgb_reg = 3'b011; end
            18'b001000001101010011: begin rgb_reg = 3'b011; end
            18'b001000001101010100: begin rgb_reg = 3'b011; end
            18'b001000001101010101: begin rgb_reg = 3'b011; end
            18'b001000001101010110: begin rgb_reg = 3'b011; end
            18'b001000001101010111: begin rgb_reg = 3'b011; end
            18'b001000001101011000: begin rgb_reg = 3'b011; end
            18'b001000001101011001: begin rgb_reg = 3'b011; end
            18'b001000001101011010: begin rgb_reg = 3'b011; end
            18'b001000001101011011: begin rgb_reg = 3'b011; end
            18'b001000001101011100: begin rgb_reg = 3'b011; end
            18'b001000001101011101: begin rgb_reg = 3'b011; end
            18'b001000001101011110: begin rgb_reg = 3'b011; end
            18'b001000001101011111: begin rgb_reg = 3'b011; end
            18'b001000001101100000: begin rgb_reg = 3'b011; end
            18'b001000001101100001: begin rgb_reg = 3'b011; end
            18'b001000001101100010: begin rgb_reg = 3'b011; end
            18'b001000001101101010: begin rgb_reg = 3'b001; end
            18'b001000001101101011: begin rgb_reg = 3'b011; end
            18'b001000001101110101: begin rgb_reg = 3'b011; end
            18'b001000001101110110: begin rgb_reg = 3'b001; end
            18'b001000010010011100: begin rgb_reg = 3'b001; end
            18'b001000010010011101: begin rgb_reg = 3'b011; end
            18'b001000010010011110: begin rgb_reg = 3'b011; end
            18'b001000010010011111: begin rgb_reg = 3'b011; end
            18'b001000010010101011: begin rgb_reg = 3'b001; end
            18'b001000010010101100: begin rgb_reg = 3'b011; end
            18'b001000010010101101: begin rgb_reg = 3'b011; end
            18'b001000010010101110: begin rgb_reg = 3'b011; end
            18'b001000010010110011: begin rgb_reg = 3'b011; end
            18'b001000010010110100: begin rgb_reg = 3'b011; end
            18'b001000010010110101: begin rgb_reg = 3'b011; end
            18'b001000010010110110: begin rgb_reg = 3'b011; end
            18'b001000010010110111: begin rgb_reg = 3'b011; end
            18'b001000010010111000: begin rgb_reg = 3'b011; end
            18'b001000010010111001: begin rgb_reg = 3'b011; end
            18'b001000010010111010: begin rgb_reg = 3'b001; end
            18'b001000010011000010: begin rgb_reg = 3'b011; end
            18'b001000010011000011: begin rgb_reg = 3'b011; end
            18'b001000010011000100: begin rgb_reg = 3'b011; end
            18'b001000010011000101: begin rgb_reg = 3'b011; end
            18'b001000010011001001: begin rgb_reg = 3'b001; end
            18'b001000010011001010: begin rgb_reg = 3'b011; end
            18'b001000010011001011: begin rgb_reg = 3'b011; end
            18'b001000010011001100: begin rgb_reg = 3'b011; end
            18'b001000010011011000: begin rgb_reg = 3'b001; end
            18'b001000010011011001: begin rgb_reg = 3'b011; end
            18'b001000010011011010: begin rgb_reg = 3'b011; end
            18'b001000010011011011: begin rgb_reg = 3'b011; end
            18'b001000010011100000: begin rgb_reg = 3'b011; end
            18'b001000010011100001: begin rgb_reg = 3'b011; end
            18'b001000010011100010: begin rgb_reg = 3'b011; end
            18'b001000010011100011: begin rgb_reg = 3'b011; end
            18'b001000010011110110: begin rgb_reg = 3'b001; end
            18'b001000010011110111: begin rgb_reg = 3'b011; end
            18'b001000010011111000: begin rgb_reg = 3'b011; end
            18'b001000010011111001: begin rgb_reg = 3'b011; end
            18'b001000010100000101: begin rgb_reg = 3'b001; end
            18'b001000010100000110: begin rgb_reg = 3'b011; end
            18'b001000010100000111: begin rgb_reg = 3'b011; end
            18'b001000010100001000: begin rgb_reg = 3'b011; end
            18'b001000010100001101: begin rgb_reg = 3'b011; end
            18'b001000010100001110: begin rgb_reg = 3'b011; end
            18'b001000010100001111: begin rgb_reg = 3'b011; end
            18'b001000010100010000: begin rgb_reg = 3'b011; end
            18'b001000010100011100: begin rgb_reg = 3'b011; end
            18'b001000010100011101: begin rgb_reg = 3'b011; end
            18'b001000010100011110: begin rgb_reg = 3'b011; end
            18'b001000010100011111: begin rgb_reg = 3'b011; end
            18'b001000010100100011: begin rgb_reg = 3'b001; end
            18'b001000010100100100: begin rgb_reg = 3'b011; end
            18'b001000010100100101: begin rgb_reg = 3'b011; end
            18'b001000010100100110: begin rgb_reg = 3'b011; end
            18'b001000010100110010: begin rgb_reg = 3'b001; end
            18'b001000010100110011: begin rgb_reg = 3'b011; end
            18'b001000010100110100: begin rgb_reg = 3'b011; end
            18'b001000010100110101: begin rgb_reg = 3'b011; end
            18'b001000010100111010: begin rgb_reg = 3'b011; end
            18'b001000010100111011: begin rgb_reg = 3'b011; end
            18'b001000010100111100: begin rgb_reg = 3'b011; end
            18'b001000010100111101: begin rgb_reg = 3'b011; end
            18'b001000010101001001: begin rgb_reg = 3'b011; end
            18'b001000010101001010: begin rgb_reg = 3'b011; end
            18'b001000010101001011: begin rgb_reg = 3'b011; end
            18'b001000010101001100: begin rgb_reg = 3'b011; end
            18'b001000010101010000: begin rgb_reg = 3'b001; end
            18'b001000010101010001: begin rgb_reg = 3'b011; end
            18'b001000010101010010: begin rgb_reg = 3'b011; end
            18'b001000010101010011: begin rgb_reg = 3'b011; end
            18'b001000010101101011: begin rgb_reg = 3'b001; end
            18'b001000010101101100: begin rgb_reg = 3'b001; end
            18'b001000010101101101: begin rgb_reg = 3'b001; end
            18'b001000010101101110: begin rgb_reg = 3'b001; end
            18'b001000010101101111: begin rgb_reg = 3'b001; end
            18'b001000010101110000: begin rgb_reg = 3'b001; end
            18'b001000010101110001: begin rgb_reg = 3'b001; end
            18'b001000010101110010: begin rgb_reg = 3'b001; end
            18'b001000010101110011: begin rgb_reg = 3'b001; end
            18'b001000010101110100: begin rgb_reg = 3'b001; end
            18'b001000010101110101: begin rgb_reg = 3'b001; end
            18'b001000011010011100: begin rgb_reg = 3'b001; end
            18'b001000011010011101: begin rgb_reg = 3'b011; end
            18'b001000011010011110: begin rgb_reg = 3'b011; end
            18'b001000011010011111: begin rgb_reg = 3'b011; end
            18'b001000011010101011: begin rgb_reg = 3'b001; end
            18'b001000011010101100: begin rgb_reg = 3'b011; end
            18'b001000011010101101: begin rgb_reg = 3'b011; end
            18'b001000011010101110: begin rgb_reg = 3'b011; end
            18'b001000011010110011: begin rgb_reg = 3'b011; end
            18'b001000011010110100: begin rgb_reg = 3'b011; end
            18'b001000011010110101: begin rgb_reg = 3'b011; end
            18'b001000011010110110: begin rgb_reg = 3'b011; end
            18'b001000011010110111: begin rgb_reg = 3'b011; end
            18'b001000011010111000: begin rgb_reg = 3'b011; end
            18'b001000011010111001: begin rgb_reg = 3'b011; end
            18'b001000011010111010: begin rgb_reg = 3'b001; end
            18'b001000011011000010: begin rgb_reg = 3'b011; end
            18'b001000011011000011: begin rgb_reg = 3'b011; end
            18'b001000011011000100: begin rgb_reg = 3'b011; end
            18'b001000011011000101: begin rgb_reg = 3'b011; end
            18'b001000011011001001: begin rgb_reg = 3'b001; end
            18'b001000011011001010: begin rgb_reg = 3'b011; end
            18'b001000011011001011: begin rgb_reg = 3'b011; end
            18'b001000011011001100: begin rgb_reg = 3'b011; end
            18'b001000011011011000: begin rgb_reg = 3'b001; end
            18'b001000011011011001: begin rgb_reg = 3'b011; end
            18'b001000011011011010: begin rgb_reg = 3'b011; end
            18'b001000011011011011: begin rgb_reg = 3'b011; end
            18'b001000011011100000: begin rgb_reg = 3'b011; end
            18'b001000011011100001: begin rgb_reg = 3'b011; end
            18'b001000011011100010: begin rgb_reg = 3'b011; end
            18'b001000011011100011: begin rgb_reg = 3'b011; end
            18'b001000011011110110: begin rgb_reg = 3'b001; end
            18'b001000011011110111: begin rgb_reg = 3'b011; end
            18'b001000011011111000: begin rgb_reg = 3'b011; end
            18'b001000011011111001: begin rgb_reg = 3'b011; end
            18'b001000011100000101: begin rgb_reg = 3'b001; end
            18'b001000011100000110: begin rgb_reg = 3'b011; end
            18'b001000011100000111: begin rgb_reg = 3'b011; end
            18'b001000011100001000: begin rgb_reg = 3'b011; end
            18'b001000011100001101: begin rgb_reg = 3'b011; end
            18'b001000011100001110: begin rgb_reg = 3'b011; end
            18'b001000011100001111: begin rgb_reg = 3'b011; end
            18'b001000011100010000: begin rgb_reg = 3'b011; end
            18'b001000011100011100: begin rgb_reg = 3'b011; end
            18'b001000011100011101: begin rgb_reg = 3'b011; end
            18'b001000011100011110: begin rgb_reg = 3'b011; end
            18'b001000011100011111: begin rgb_reg = 3'b011; end
            18'b001000011100100011: begin rgb_reg = 3'b001; end
            18'b001000011100100100: begin rgb_reg = 3'b011; end
            18'b001000011100100101: begin rgb_reg = 3'b011; end
            18'b001000011100100110: begin rgb_reg = 3'b011; end
            18'b001000011100110010: begin rgb_reg = 3'b001; end
            18'b001000011100110011: begin rgb_reg = 3'b011; end
            18'b001000011100110100: begin rgb_reg = 3'b011; end
            18'b001000011100110101: begin rgb_reg = 3'b011; end
            18'b001000011100111010: begin rgb_reg = 3'b011; end
            18'b001000011100111011: begin rgb_reg = 3'b011; end
            18'b001000011100111100: begin rgb_reg = 3'b011; end
            18'b001000011100111101: begin rgb_reg = 3'b011; end
            18'b001000011101001001: begin rgb_reg = 3'b011; end
            18'b001000011101001010: begin rgb_reg = 3'b011; end
            18'b001000011101001011: begin rgb_reg = 3'b011; end
            18'b001000011101001100: begin rgb_reg = 3'b011; end
            18'b001000011101010000: begin rgb_reg = 3'b001; end
            18'b001000011101010001: begin rgb_reg = 3'b011; end
            18'b001000011101010010: begin rgb_reg = 3'b011; end
            18'b001000011101010011: begin rgb_reg = 3'b011; end
            18'b001000011101101100: begin rgb_reg = 3'b001; end
            18'b001000011101101101: begin rgb_reg = 3'b011; end
            18'b001000011101101110: begin rgb_reg = 3'b011; end
            18'b001000011101101111: begin rgb_reg = 3'b011; end
            18'b001000011101110000: begin rgb_reg = 3'b011; end
            18'b001000011101110001: begin rgb_reg = 3'b011; end
            18'b001000011101110010: begin rgb_reg = 3'b011; end
            18'b001000011101110011: begin rgb_reg = 3'b011; end
            18'b001000011101110100: begin rgb_reg = 3'b011; end
            18'b001000100010011100: begin rgb_reg = 3'b001; end
            18'b001000100010011101: begin rgb_reg = 3'b011; end
            18'b001000100010011110: begin rgb_reg = 3'b011; end
            18'b001000100010011111: begin rgb_reg = 3'b011; end
            18'b001000100010101011: begin rgb_reg = 3'b001; end
            18'b001000100010101100: begin rgb_reg = 3'b011; end
            18'b001000100010101101: begin rgb_reg = 3'b011; end
            18'b001000100010101110: begin rgb_reg = 3'b011; end
            18'b001000100010110011: begin rgb_reg = 3'b011; end
            18'b001000100010110100: begin rgb_reg = 3'b011; end
            18'b001000100010110101: begin rgb_reg = 3'b011; end
            18'b001000100010110110: begin rgb_reg = 3'b011; end
            18'b001000100010110111: begin rgb_reg = 3'b011; end
            18'b001000100010111000: begin rgb_reg = 3'b011; end
            18'b001000100010111001: begin rgb_reg = 3'b011; end
            18'b001000100010111010: begin rgb_reg = 3'b001; end
            18'b001000100011000010: begin rgb_reg = 3'b011; end
            18'b001000100011000011: begin rgb_reg = 3'b011; end
            18'b001000100011000100: begin rgb_reg = 3'b011; end
            18'b001000100011000101: begin rgb_reg = 3'b011; end
            18'b001000100011001001: begin rgb_reg = 3'b001; end
            18'b001000100011001010: begin rgb_reg = 3'b011; end
            18'b001000100011001011: begin rgb_reg = 3'b011; end
            18'b001000100011001100: begin rgb_reg = 3'b011; end
            18'b001000100011011000: begin rgb_reg = 3'b001; end
            18'b001000100011011001: begin rgb_reg = 3'b011; end
            18'b001000100011011010: begin rgb_reg = 3'b011; end
            18'b001000100011011011: begin rgb_reg = 3'b011; end
            18'b001000100011100000: begin rgb_reg = 3'b011; end
            18'b001000100011100001: begin rgb_reg = 3'b011; end
            18'b001000100011100010: begin rgb_reg = 3'b011; end
            18'b001000100011100011: begin rgb_reg = 3'b011; end
            18'b001000100011110110: begin rgb_reg = 3'b001; end
            18'b001000100011110111: begin rgb_reg = 3'b011; end
            18'b001000100011111000: begin rgb_reg = 3'b011; end
            18'b001000100011111001: begin rgb_reg = 3'b011; end
            18'b001000100100000101: begin rgb_reg = 3'b001; end
            18'b001000100100000110: begin rgb_reg = 3'b011; end
            18'b001000100100000111: begin rgb_reg = 3'b011; end
            18'b001000100100001000: begin rgb_reg = 3'b011; end
            18'b001000100100001101: begin rgb_reg = 3'b011; end
            18'b001000100100001110: begin rgb_reg = 3'b011; end
            18'b001000100100001111: begin rgb_reg = 3'b011; end
            18'b001000100100010000: begin rgb_reg = 3'b011; end
            18'b001000100100011100: begin rgb_reg = 3'b011; end
            18'b001000100100011101: begin rgb_reg = 3'b011; end
            18'b001000100100011110: begin rgb_reg = 3'b011; end
            18'b001000100100011111: begin rgb_reg = 3'b011; end
            18'b001000100100100011: begin rgb_reg = 3'b001; end
            18'b001000100100100100: begin rgb_reg = 3'b011; end
            18'b001000100100100101: begin rgb_reg = 3'b011; end
            18'b001000100100100110: begin rgb_reg = 3'b011; end
            18'b001000100100110010: begin rgb_reg = 3'b001; end
            18'b001000100100110011: begin rgb_reg = 3'b011; end
            18'b001000100100110100: begin rgb_reg = 3'b011; end
            18'b001000100100110101: begin rgb_reg = 3'b011; end
            18'b001000100100111010: begin rgb_reg = 3'b011; end
            18'b001000100100111011: begin rgb_reg = 3'b011; end
            18'b001000100100111100: begin rgb_reg = 3'b011; end
            18'b001000100100111101: begin rgb_reg = 3'b011; end
            18'b001000100101001001: begin rgb_reg = 3'b011; end
            18'b001000100101001010: begin rgb_reg = 3'b011; end
            18'b001000100101001011: begin rgb_reg = 3'b011; end
            18'b001000100101001100: begin rgb_reg = 3'b011; end
            18'b001000100101010000: begin rgb_reg = 3'b001; end
            18'b001000100101010001: begin rgb_reg = 3'b011; end
            18'b001000100101010010: begin rgb_reg = 3'b011; end
            18'b001000100101010011: begin rgb_reg = 3'b011; end
            18'b001000101010011100: begin rgb_reg = 3'b001; end
            18'b001000101010011101: begin rgb_reg = 3'b011; end
            18'b001000101010011110: begin rgb_reg = 3'b011; end
            18'b001000101010011111: begin rgb_reg = 3'b011; end
            18'b001000101010101011: begin rgb_reg = 3'b001; end
            18'b001000101010101100: begin rgb_reg = 3'b011; end
            18'b001000101010101101: begin rgb_reg = 3'b011; end
            18'b001000101010101110: begin rgb_reg = 3'b011; end
            18'b001000101010110011: begin rgb_reg = 3'b011; end
            18'b001000101010110100: begin rgb_reg = 3'b011; end
            18'b001000101010110101: begin rgb_reg = 3'b011; end
            18'b001000101010110110: begin rgb_reg = 3'b011; end
            18'b001000101010110111: begin rgb_reg = 3'b001; end
            18'b001000101010111000: begin rgb_reg = 3'b001; end
            18'b001000101010111001: begin rgb_reg = 3'b001; end
            18'b001000101010111010: begin rgb_reg = 3'b001; end
            18'b001000101010111011: begin rgb_reg = 3'b001; end
            18'b001000101010111100: begin rgb_reg = 3'b001; end
            18'b001000101010111101: begin rgb_reg = 3'b001; end
            18'b001000101011000010: begin rgb_reg = 3'b011; end
            18'b001000101011000011: begin rgb_reg = 3'b011; end
            18'b001000101011000100: begin rgb_reg = 3'b011; end
            18'b001000101011000101: begin rgb_reg = 3'b011; end
            18'b001000101011001001: begin rgb_reg = 3'b001; end
            18'b001000101011001010: begin rgb_reg = 3'b011; end
            18'b001000101011001011: begin rgb_reg = 3'b011; end
            18'b001000101011001100: begin rgb_reg = 3'b011; end
            18'b001000101011011000: begin rgb_reg = 3'b001; end
            18'b001000101011011001: begin rgb_reg = 3'b011; end
            18'b001000101011011010: begin rgb_reg = 3'b011; end
            18'b001000101011011011: begin rgb_reg = 3'b011; end
            18'b001000101011100000: begin rgb_reg = 3'b011; end
            18'b001000101011100001: begin rgb_reg = 3'b011; end
            18'b001000101011100010: begin rgb_reg = 3'b011; end
            18'b001000101011100011: begin rgb_reg = 3'b011; end
            18'b001000101011100100: begin rgb_reg = 3'b001; end
            18'b001000101011100101: begin rgb_reg = 3'b001; end
            18'b001000101011100110: begin rgb_reg = 3'b001; end
            18'b001000101011100111: begin rgb_reg = 3'b001; end
            18'b001000101011101000: begin rgb_reg = 3'b001; end
            18'b001000101011101001: begin rgb_reg = 3'b001; end
            18'b001000101011101010: begin rgb_reg = 3'b001; end
            18'b001000101011110110: begin rgb_reg = 3'b001; end
            18'b001000101011110111: begin rgb_reg = 3'b011; end
            18'b001000101011111000: begin rgb_reg = 3'b011; end
            18'b001000101011111001: begin rgb_reg = 3'b011; end
            18'b001000101011111010: begin rgb_reg = 3'b001; end
            18'b001000101011111011: begin rgb_reg = 3'b001; end
            18'b001000101011111100: begin rgb_reg = 3'b001; end
            18'b001000101011111101: begin rgb_reg = 3'b001; end
            18'b001000101011111110: begin rgb_reg = 3'b001; end
            18'b001000101011111111: begin rgb_reg = 3'b001; end
            18'b001000101100000000: begin rgb_reg = 3'b001; end
            18'b001000101100000001: begin rgb_reg = 3'b001; end
            18'b001000101100000010: begin rgb_reg = 3'b001; end
            18'b001000101100000011: begin rgb_reg = 3'b001; end
            18'b001000101100000100: begin rgb_reg = 3'b001; end
            18'b001000101100000101: begin rgb_reg = 3'b001; end
            18'b001000101100000110: begin rgb_reg = 3'b001; end
            18'b001000101100000111: begin rgb_reg = 3'b001; end
            18'b001000101100001000: begin rgb_reg = 3'b001; end
            18'b001000101100001101: begin rgb_reg = 3'b011; end
            18'b001000101100001110: begin rgb_reg = 3'b011; end
            18'b001000101100001111: begin rgb_reg = 3'b011; end
            18'b001000101100010000: begin rgb_reg = 3'b011; end
            18'b001000101100011100: begin rgb_reg = 3'b011; end
            18'b001000101100011101: begin rgb_reg = 3'b011; end
            18'b001000101100011110: begin rgb_reg = 3'b011; end
            18'b001000101100011111: begin rgb_reg = 3'b011; end
            18'b001000101100100011: begin rgb_reg = 3'b001; end
            18'b001000101100100100: begin rgb_reg = 3'b011; end
            18'b001000101100100101: begin rgb_reg = 3'b011; end
            18'b001000101100100110: begin rgb_reg = 3'b011; end
            18'b001000101100100111: begin rgb_reg = 3'b001; end
            18'b001000101100101000: begin rgb_reg = 3'b001; end
            18'b001000101100101001: begin rgb_reg = 3'b001; end
            18'b001000101100101010: begin rgb_reg = 3'b001; end
            18'b001000101100101011: begin rgb_reg = 3'b001; end
            18'b001000101100101100: begin rgb_reg = 3'b001; end
            18'b001000101100101101: begin rgb_reg = 3'b001; end
            18'b001000101100101110: begin rgb_reg = 3'b001; end
            18'b001000101100101111: begin rgb_reg = 3'b001; end
            18'b001000101100110000: begin rgb_reg = 3'b001; end
            18'b001000101100110001: begin rgb_reg = 3'b001; end
            18'b001000101100110010: begin rgb_reg = 3'b011; end
            18'b001000101100110011: begin rgb_reg = 3'b011; end
            18'b001000101100110100: begin rgb_reg = 3'b011; end
            18'b001000101100110101: begin rgb_reg = 3'b011; end
            18'b001000101100111010: begin rgb_reg = 3'b011; end
            18'b001000101100111011: begin rgb_reg = 3'b011; end
            18'b001000101100111100: begin rgb_reg = 3'b011; end
            18'b001000101100111101: begin rgb_reg = 3'b011; end
            18'b001000101100111110: begin rgb_reg = 3'b001; end
            18'b001000101100111111: begin rgb_reg = 3'b001; end
            18'b001000101101000000: begin rgb_reg = 3'b001; end
            18'b001000101101000001: begin rgb_reg = 3'b001; end
            18'b001000101101000010: begin rgb_reg = 3'b001; end
            18'b001000101101000011: begin rgb_reg = 3'b001; end
            18'b001000101101000100: begin rgb_reg = 3'b001; end
            18'b001000101101000101: begin rgb_reg = 3'b001; end
            18'b001000101101000110: begin rgb_reg = 3'b001; end
            18'b001000101101000111: begin rgb_reg = 3'b001; end
            18'b001000101101001000: begin rgb_reg = 3'b001; end
            18'b001000101101001001: begin rgb_reg = 3'b001; end
            18'b001000101101001010: begin rgb_reg = 3'b001; end
            18'b001000101101001011: begin rgb_reg = 3'b001; end
            18'b001000101101001100: begin rgb_reg = 3'b001; end
            18'b001000101101010000: begin rgb_reg = 3'b001; end
            18'b001000101101010001: begin rgb_reg = 3'b011; end
            18'b001000101101010010: begin rgb_reg = 3'b011; end
            18'b001000101101010011: begin rgb_reg = 3'b011; end
            18'b001000101101010100: begin rgb_reg = 3'b001; end
            18'b001000101101010101: begin rgb_reg = 3'b001; end
            18'b001000101101010110: begin rgb_reg = 3'b001; end
            18'b001000101101010111: begin rgb_reg = 3'b001; end
            18'b001000101101011000: begin rgb_reg = 3'b001; end
            18'b001000101101011001: begin rgb_reg = 3'b001; end
            18'b001000101101011010: begin rgb_reg = 3'b001; end
            18'b001000101101011011: begin rgb_reg = 3'b001; end
            18'b001000110010011100: begin rgb_reg = 3'b001; end
            18'b001000110010011101: begin rgb_reg = 3'b011; end
            18'b001000110010011110: begin rgb_reg = 3'b011; end
            18'b001000110010011111: begin rgb_reg = 3'b011; end
            18'b001000110010101011: begin rgb_reg = 3'b001; end
            18'b001000110010101100: begin rgb_reg = 3'b011; end
            18'b001000110010101101: begin rgb_reg = 3'b011; end
            18'b001000110010101110: begin rgb_reg = 3'b011; end
            18'b001000110010110011: begin rgb_reg = 3'b011; end
            18'b001000110010110100: begin rgb_reg = 3'b011; end
            18'b001000110010110101: begin rgb_reg = 3'b011; end
            18'b001000110010110110: begin rgb_reg = 3'b011; end
            18'b001000110010111010: begin rgb_reg = 3'b001; end
            18'b001000110010111011: begin rgb_reg = 3'b011; end
            18'b001000110010111100: begin rgb_reg = 3'b011; end
            18'b001000110010111101: begin rgb_reg = 3'b011; end
            18'b001000110011000010: begin rgb_reg = 3'b011; end
            18'b001000110011000011: begin rgb_reg = 3'b011; end
            18'b001000110011000100: begin rgb_reg = 3'b011; end
            18'b001000110011000101: begin rgb_reg = 3'b011; end
            18'b001000110011001001: begin rgb_reg = 3'b001; end
            18'b001000110011001010: begin rgb_reg = 3'b011; end
            18'b001000110011001011: begin rgb_reg = 3'b011; end
            18'b001000110011001100: begin rgb_reg = 3'b011; end
            18'b001000110011011000: begin rgb_reg = 3'b001; end
            18'b001000110011011001: begin rgb_reg = 3'b011; end
            18'b001000110011011010: begin rgb_reg = 3'b011; end
            18'b001000110011011011: begin rgb_reg = 3'b011; end
            18'b001000110011100000: begin rgb_reg = 3'b011; end
            18'b001000110011100001: begin rgb_reg = 3'b011; end
            18'b001000110011100010: begin rgb_reg = 3'b011; end
            18'b001000110011100011: begin rgb_reg = 3'b011; end
            18'b001000110011100100: begin rgb_reg = 3'b011; end
            18'b001000110011100101: begin rgb_reg = 3'b011; end
            18'b001000110011100110: begin rgb_reg = 3'b011; end
            18'b001000110011100111: begin rgb_reg = 3'b011; end
            18'b001000110011101000: begin rgb_reg = 3'b011; end
            18'b001000110011101001: begin rgb_reg = 3'b011; end
            18'b001000110011101010: begin rgb_reg = 3'b011; end
            18'b001000110011110110: begin rgb_reg = 3'b001; end
            18'b001000110011110111: begin rgb_reg = 3'b011; end
            18'b001000110011111000: begin rgb_reg = 3'b011; end
            18'b001000110011111001: begin rgb_reg = 3'b011; end
            18'b001000110011111010: begin rgb_reg = 3'b011; end
            18'b001000110011111011: begin rgb_reg = 3'b011; end
            18'b001000110011111100: begin rgb_reg = 3'b011; end
            18'b001000110011111101: begin rgb_reg = 3'b011; end
            18'b001000110011111110: begin rgb_reg = 3'b011; end
            18'b001000110011111111: begin rgb_reg = 3'b011; end
            18'b001000110100000000: begin rgb_reg = 3'b011; end
            18'b001000110100000001: begin rgb_reg = 3'b011; end
            18'b001000110100000010: begin rgb_reg = 3'b011; end
            18'b001000110100000011: begin rgb_reg = 3'b011; end
            18'b001000110100000100: begin rgb_reg = 3'b011; end
            18'b001000110100000101: begin rgb_reg = 3'b001; end
            18'b001000110100001101: begin rgb_reg = 3'b011; end
            18'b001000110100001110: begin rgb_reg = 3'b011; end
            18'b001000110100001111: begin rgb_reg = 3'b011; end
            18'b001000110100010000: begin rgb_reg = 3'b011; end
            18'b001000110100011100: begin rgb_reg = 3'b011; end
            18'b001000110100011101: begin rgb_reg = 3'b011; end
            18'b001000110100011110: begin rgb_reg = 3'b011; end
            18'b001000110100011111: begin rgb_reg = 3'b011; end
            18'b001000110100100011: begin rgb_reg = 3'b001; end
            18'b001000110100100100: begin rgb_reg = 3'b011; end
            18'b001000110100100101: begin rgb_reg = 3'b011; end
            18'b001000110100100110: begin rgb_reg = 3'b011; end
            18'b001000110100100111: begin rgb_reg = 3'b011; end
            18'b001000110100101000: begin rgb_reg = 3'b011; end
            18'b001000110100101001: begin rgb_reg = 3'b011; end
            18'b001000110100101010: begin rgb_reg = 3'b011; end
            18'b001000110100101011: begin rgb_reg = 3'b011; end
            18'b001000110100101100: begin rgb_reg = 3'b011; end
            18'b001000110100101101: begin rgb_reg = 3'b011; end
            18'b001000110100101110: begin rgb_reg = 3'b011; end
            18'b001000110100101111: begin rgb_reg = 3'b011; end
            18'b001000110100110000: begin rgb_reg = 3'b011; end
            18'b001000110100110001: begin rgb_reg = 3'b011; end
            18'b001000110100110010: begin rgb_reg = 3'b011; end
            18'b001000110100110011: begin rgb_reg = 3'b011; end
            18'b001000110100110100: begin rgb_reg = 3'b011; end
            18'b001000110100110101: begin rgb_reg = 3'b011; end
            18'b001000110100111010: begin rgb_reg = 3'b011; end
            18'b001000110100111011: begin rgb_reg = 3'b011; end
            18'b001000110100111100: begin rgb_reg = 3'b011; end
            18'b001000110100111101: begin rgb_reg = 3'b011; end
            18'b001000110100111110: begin rgb_reg = 3'b011; end
            18'b001000110100111111: begin rgb_reg = 3'b011; end
            18'b001000110101000000: begin rgb_reg = 3'b011; end
            18'b001000110101000001: begin rgb_reg = 3'b011; end
            18'b001000110101000010: begin rgb_reg = 3'b011; end
            18'b001000110101000011: begin rgb_reg = 3'b011; end
            18'b001000110101000100: begin rgb_reg = 3'b011; end
            18'b001000110101000101: begin rgb_reg = 3'b011; end
            18'b001000110101000110: begin rgb_reg = 3'b011; end
            18'b001000110101000111: begin rgb_reg = 3'b011; end
            18'b001000110101001000: begin rgb_reg = 3'b011; end
            18'b001000110101010000: begin rgb_reg = 3'b001; end
            18'b001000110101010001: begin rgb_reg = 3'b011; end
            18'b001000110101010010: begin rgb_reg = 3'b011; end
            18'b001000110101010011: begin rgb_reg = 3'b011; end
            18'b001000110101010100: begin rgb_reg = 3'b011; end
            18'b001000110101010101: begin rgb_reg = 3'b011; end
            18'b001000110101010110: begin rgb_reg = 3'b011; end
            18'b001000110101010111: begin rgb_reg = 3'b011; end
            18'b001000110101011000: begin rgb_reg = 3'b011; end
            18'b001000110101011001: begin rgb_reg = 3'b011; end
            18'b001000110101011010: begin rgb_reg = 3'b011; end
            18'b001000110101011011: begin rgb_reg = 3'b011; end
            18'b001000111010011100: begin rgb_reg = 3'b001; end
            18'b001000111010011101: begin rgb_reg = 3'b011; end
            18'b001000111010011110: begin rgb_reg = 3'b011; end
            18'b001000111010011111: begin rgb_reg = 3'b011; end
            18'b001000111010101011: begin rgb_reg = 3'b001; end
            18'b001000111010101100: begin rgb_reg = 3'b011; end
            18'b001000111010101101: begin rgb_reg = 3'b011; end
            18'b001000111010101110: begin rgb_reg = 3'b011; end
            18'b001000111010110011: begin rgb_reg = 3'b011; end
            18'b001000111010110100: begin rgb_reg = 3'b011; end
            18'b001000111010110101: begin rgb_reg = 3'b011; end
            18'b001000111010110110: begin rgb_reg = 3'b011; end
            18'b001000111010111010: begin rgb_reg = 3'b001; end
            18'b001000111010111011: begin rgb_reg = 3'b011; end
            18'b001000111010111100: begin rgb_reg = 3'b011; end
            18'b001000111010111101: begin rgb_reg = 3'b011; end
            18'b001000111011000010: begin rgb_reg = 3'b011; end
            18'b001000111011000011: begin rgb_reg = 3'b011; end
            18'b001000111011000100: begin rgb_reg = 3'b011; end
            18'b001000111011000101: begin rgb_reg = 3'b011; end
            18'b001000111011001001: begin rgb_reg = 3'b001; end
            18'b001000111011001010: begin rgb_reg = 3'b011; end
            18'b001000111011001011: begin rgb_reg = 3'b011; end
            18'b001000111011001100: begin rgb_reg = 3'b011; end
            18'b001000111011011000: begin rgb_reg = 3'b001; end
            18'b001000111011011001: begin rgb_reg = 3'b011; end
            18'b001000111011011010: begin rgb_reg = 3'b011; end
            18'b001000111011011011: begin rgb_reg = 3'b011; end
            18'b001000111011100000: begin rgb_reg = 3'b011; end
            18'b001000111011100001: begin rgb_reg = 3'b011; end
            18'b001000111011100010: begin rgb_reg = 3'b011; end
            18'b001000111011100011: begin rgb_reg = 3'b011; end
            18'b001000111011100100: begin rgb_reg = 3'b011; end
            18'b001000111011100101: begin rgb_reg = 3'b011; end
            18'b001000111011100110: begin rgb_reg = 3'b011; end
            18'b001000111011100111: begin rgb_reg = 3'b011; end
            18'b001000111011101000: begin rgb_reg = 3'b011; end
            18'b001000111011101001: begin rgb_reg = 3'b011; end
            18'b001000111011101010: begin rgb_reg = 3'b011; end
            18'b001000111011110110: begin rgb_reg = 3'b001; end
            18'b001000111011110111: begin rgb_reg = 3'b011; end
            18'b001000111011111000: begin rgb_reg = 3'b011; end
            18'b001000111011111001: begin rgb_reg = 3'b011; end
            18'b001000111011111010: begin rgb_reg = 3'b011; end
            18'b001000111011111011: begin rgb_reg = 3'b011; end
            18'b001000111011111100: begin rgb_reg = 3'b011; end
            18'b001000111011111101: begin rgb_reg = 3'b011; end
            18'b001000111011111110: begin rgb_reg = 3'b011; end
            18'b001000111011111111: begin rgb_reg = 3'b011; end
            18'b001000111100000000: begin rgb_reg = 3'b011; end
            18'b001000111100000001: begin rgb_reg = 3'b011; end
            18'b001000111100000010: begin rgb_reg = 3'b011; end
            18'b001000111100000011: begin rgb_reg = 3'b011; end
            18'b001000111100000100: begin rgb_reg = 3'b011; end
            18'b001000111100000101: begin rgb_reg = 3'b001; end
            18'b001000111100001101: begin rgb_reg = 3'b011; end
            18'b001000111100001110: begin rgb_reg = 3'b011; end
            18'b001000111100001111: begin rgb_reg = 3'b011; end
            18'b001000111100010000: begin rgb_reg = 3'b011; end
            18'b001000111100011100: begin rgb_reg = 3'b011; end
            18'b001000111100011101: begin rgb_reg = 3'b011; end
            18'b001000111100011110: begin rgb_reg = 3'b011; end
            18'b001000111100011111: begin rgb_reg = 3'b011; end
            18'b001000111100100011: begin rgb_reg = 3'b001; end
            18'b001000111100100100: begin rgb_reg = 3'b011; end
            18'b001000111100100101: begin rgb_reg = 3'b011; end
            18'b001000111100100110: begin rgb_reg = 3'b011; end
            18'b001000111100100111: begin rgb_reg = 3'b011; end
            18'b001000111100101000: begin rgb_reg = 3'b011; end
            18'b001000111100101001: begin rgb_reg = 3'b011; end
            18'b001000111100101010: begin rgb_reg = 3'b011; end
            18'b001000111100101011: begin rgb_reg = 3'b011; end
            18'b001000111100101100: begin rgb_reg = 3'b011; end
            18'b001000111100101101: begin rgb_reg = 3'b011; end
            18'b001000111100101110: begin rgb_reg = 3'b011; end
            18'b001000111100101111: begin rgb_reg = 3'b011; end
            18'b001000111100110000: begin rgb_reg = 3'b011; end
            18'b001000111100110001: begin rgb_reg = 3'b011; end
            18'b001000111100110010: begin rgb_reg = 3'b011; end
            18'b001000111100110011: begin rgb_reg = 3'b011; end
            18'b001000111100110100: begin rgb_reg = 3'b011; end
            18'b001000111100110101: begin rgb_reg = 3'b011; end
            18'b001000111100111010: begin rgb_reg = 3'b011; end
            18'b001000111100111011: begin rgb_reg = 3'b011; end
            18'b001000111100111100: begin rgb_reg = 3'b011; end
            18'b001000111100111101: begin rgb_reg = 3'b011; end
            18'b001000111100111110: begin rgb_reg = 3'b011; end
            18'b001000111100111111: begin rgb_reg = 3'b011; end
            18'b001000111101000000: begin rgb_reg = 3'b011; end
            18'b001000111101000001: begin rgb_reg = 3'b011; end
            18'b001000111101000010: begin rgb_reg = 3'b011; end
            18'b001000111101000011: begin rgb_reg = 3'b011; end
            18'b001000111101000100: begin rgb_reg = 3'b011; end
            18'b001000111101000101: begin rgb_reg = 3'b011; end
            18'b001000111101000110: begin rgb_reg = 3'b011; end
            18'b001000111101000111: begin rgb_reg = 3'b011; end
            18'b001000111101001000: begin rgb_reg = 3'b011; end
            18'b001000111101010000: begin rgb_reg = 3'b001; end
            18'b001000111101010001: begin rgb_reg = 3'b011; end
            18'b001000111101010010: begin rgb_reg = 3'b011; end
            18'b001000111101010011: begin rgb_reg = 3'b011; end
            18'b001000111101010100: begin rgb_reg = 3'b011; end
            18'b001000111101010101: begin rgb_reg = 3'b011; end
            18'b001000111101010110: begin rgb_reg = 3'b011; end
            18'b001000111101010111: begin rgb_reg = 3'b011; end
            18'b001000111101011000: begin rgb_reg = 3'b011; end
            18'b001000111101011001: begin rgb_reg = 3'b011; end
            18'b001000111101011010: begin rgb_reg = 3'b011; end
            18'b001000111101011011: begin rgb_reg = 3'b011; end
            18'b001001000010011100: begin rgb_reg = 3'b001; end
            18'b001001000010011101: begin rgb_reg = 3'b011; end
            18'b001001000010011110: begin rgb_reg = 3'b011; end
            18'b001001000010011111: begin rgb_reg = 3'b011; end
            18'b001001000010101011: begin rgb_reg = 3'b001; end
            18'b001001000010101100: begin rgb_reg = 3'b011; end
            18'b001001000010101101: begin rgb_reg = 3'b011; end
            18'b001001000010101110: begin rgb_reg = 3'b011; end
            18'b001001000010110011: begin rgb_reg = 3'b011; end
            18'b001001000010110100: begin rgb_reg = 3'b011; end
            18'b001001000010110101: begin rgb_reg = 3'b011; end
            18'b001001000010110110: begin rgb_reg = 3'b011; end
            18'b001001000010111010: begin rgb_reg = 3'b001; end
            18'b001001000010111011: begin rgb_reg = 3'b011; end
            18'b001001000010111100: begin rgb_reg = 3'b011; end
            18'b001001000010111101: begin rgb_reg = 3'b011; end
            18'b001001000011000010: begin rgb_reg = 3'b011; end
            18'b001001000011000011: begin rgb_reg = 3'b011; end
            18'b001001000011000100: begin rgb_reg = 3'b011; end
            18'b001001000011000101: begin rgb_reg = 3'b011; end
            18'b001001000011001001: begin rgb_reg = 3'b001; end
            18'b001001000011001010: begin rgb_reg = 3'b011; end
            18'b001001000011001011: begin rgb_reg = 3'b011; end
            18'b001001000011001100: begin rgb_reg = 3'b011; end
            18'b001001000011011000: begin rgb_reg = 3'b001; end
            18'b001001000011011001: begin rgb_reg = 3'b011; end
            18'b001001000011011010: begin rgb_reg = 3'b011; end
            18'b001001000011011011: begin rgb_reg = 3'b011; end
            18'b001001000011100000: begin rgb_reg = 3'b011; end
            18'b001001000011100001: begin rgb_reg = 3'b011; end
            18'b001001000011100010: begin rgb_reg = 3'b011; end
            18'b001001000011100011: begin rgb_reg = 3'b011; end
            18'b001001000011100100: begin rgb_reg = 3'b011; end
            18'b001001000011100101: begin rgb_reg = 3'b011; end
            18'b001001000011100110: begin rgb_reg = 3'b011; end
            18'b001001000011100111: begin rgb_reg = 3'b011; end
            18'b001001000011101000: begin rgb_reg = 3'b011; end
            18'b001001000011101001: begin rgb_reg = 3'b011; end
            18'b001001000011101010: begin rgb_reg = 3'b011; end
            18'b001001000011110110: begin rgb_reg = 3'b001; end
            18'b001001000011110111: begin rgb_reg = 3'b011; end
            18'b001001000011111000: begin rgb_reg = 3'b011; end
            18'b001001000011111001: begin rgb_reg = 3'b011; end
            18'b001001000011111010: begin rgb_reg = 3'b011; end
            18'b001001000011111011: begin rgb_reg = 3'b011; end
            18'b001001000011111100: begin rgb_reg = 3'b011; end
            18'b001001000011111101: begin rgb_reg = 3'b011; end
            18'b001001000011111110: begin rgb_reg = 3'b011; end
            18'b001001000011111111: begin rgb_reg = 3'b011; end
            18'b001001000100000000: begin rgb_reg = 3'b011; end
            18'b001001000100000001: begin rgb_reg = 3'b011; end
            18'b001001000100000010: begin rgb_reg = 3'b011; end
            18'b001001000100000011: begin rgb_reg = 3'b011; end
            18'b001001000100000100: begin rgb_reg = 3'b011; end
            18'b001001000100000101: begin rgb_reg = 3'b001; end
            18'b001001000100001101: begin rgb_reg = 3'b011; end
            18'b001001000100001110: begin rgb_reg = 3'b011; end
            18'b001001000100001111: begin rgb_reg = 3'b011; end
            18'b001001000100010000: begin rgb_reg = 3'b011; end
            18'b001001000100011100: begin rgb_reg = 3'b011; end
            18'b001001000100011101: begin rgb_reg = 3'b011; end
            18'b001001000100011110: begin rgb_reg = 3'b011; end
            18'b001001000100011111: begin rgb_reg = 3'b011; end
            18'b001001000100100011: begin rgb_reg = 3'b001; end
            18'b001001000100100100: begin rgb_reg = 3'b011; end
            18'b001001000100100101: begin rgb_reg = 3'b011; end
            18'b001001000100100110: begin rgb_reg = 3'b011; end
            18'b001001000100100111: begin rgb_reg = 3'b011; end
            18'b001001000100101000: begin rgb_reg = 3'b011; end
            18'b001001000100101001: begin rgb_reg = 3'b011; end
            18'b001001000100101010: begin rgb_reg = 3'b011; end
            18'b001001000100101011: begin rgb_reg = 3'b011; end
            18'b001001000100101100: begin rgb_reg = 3'b011; end
            18'b001001000100101101: begin rgb_reg = 3'b011; end
            18'b001001000100101110: begin rgb_reg = 3'b011; end
            18'b001001000100101111: begin rgb_reg = 3'b011; end
            18'b001001000100110000: begin rgb_reg = 3'b011; end
            18'b001001000100110001: begin rgb_reg = 3'b011; end
            18'b001001000100110010: begin rgb_reg = 3'b011; end
            18'b001001000100110011: begin rgb_reg = 3'b011; end
            18'b001001000100110100: begin rgb_reg = 3'b011; end
            18'b001001000100110101: begin rgb_reg = 3'b011; end
            18'b001001000100111010: begin rgb_reg = 3'b011; end
            18'b001001000100111011: begin rgb_reg = 3'b011; end
            18'b001001000100111100: begin rgb_reg = 3'b011; end
            18'b001001000100111101: begin rgb_reg = 3'b011; end
            18'b001001000100111110: begin rgb_reg = 3'b011; end
            18'b001001000100111111: begin rgb_reg = 3'b011; end
            18'b001001000101000000: begin rgb_reg = 3'b011; end
            18'b001001000101000001: begin rgb_reg = 3'b011; end
            18'b001001000101000010: begin rgb_reg = 3'b011; end
            18'b001001000101000011: begin rgb_reg = 3'b011; end
            18'b001001000101000100: begin rgb_reg = 3'b011; end
            18'b001001000101000101: begin rgb_reg = 3'b011; end
            18'b001001000101000110: begin rgb_reg = 3'b011; end
            18'b001001000101000111: begin rgb_reg = 3'b011; end
            18'b001001000101001000: begin rgb_reg = 3'b011; end
            18'b001001000101010000: begin rgb_reg = 3'b001; end
            18'b001001000101010001: begin rgb_reg = 3'b011; end
            18'b001001000101010010: begin rgb_reg = 3'b011; end
            18'b001001000101010011: begin rgb_reg = 3'b011; end
            18'b001001000101010100: begin rgb_reg = 3'b011; end
            18'b001001000101010101: begin rgb_reg = 3'b011; end
            18'b001001000101010110: begin rgb_reg = 3'b011; end
            18'b001001000101010111: begin rgb_reg = 3'b011; end
            18'b001001000101011000: begin rgb_reg = 3'b011; end
            18'b001001000101011001: begin rgb_reg = 3'b011; end
            18'b001001000101011010: begin rgb_reg = 3'b011; end
            18'b001001000101011011: begin rgb_reg = 3'b011; end
            18'b001001001010011100: begin rgb_reg = 3'b001; end
            18'b001001001010011101: begin rgb_reg = 3'b011; end
            18'b001001001010011110: begin rgb_reg = 3'b011; end
            18'b001001001010011111: begin rgb_reg = 3'b011; end
            18'b001001001010101011: begin rgb_reg = 3'b001; end
            18'b001001001010101100: begin rgb_reg = 3'b011; end
            18'b001001001010101101: begin rgb_reg = 3'b011; end
            18'b001001001010101110: begin rgb_reg = 3'b011; end
            18'b001001001010110011: begin rgb_reg = 3'b011; end
            18'b001001001010110100: begin rgb_reg = 3'b011; end
            18'b001001001010110101: begin rgb_reg = 3'b011; end
            18'b001001001010110110: begin rgb_reg = 3'b011; end
            18'b001001001010111110: begin rgb_reg = 3'b001; end
            18'b001001001010111111: begin rgb_reg = 3'b011; end
            18'b001001001011000000: begin rgb_reg = 3'b011; end
            18'b001001001011000001: begin rgb_reg = 3'b011; end
            18'b001001001011000010: begin rgb_reg = 3'b011; end
            18'b001001001011000011: begin rgb_reg = 3'b011; end
            18'b001001001011000100: begin rgb_reg = 3'b011; end
            18'b001001001011000101: begin rgb_reg = 3'b011; end
            18'b001001001011001001: begin rgb_reg = 3'b001; end
            18'b001001001011001010: begin rgb_reg = 3'b011; end
            18'b001001001011001011: begin rgb_reg = 3'b011; end
            18'b001001001011001100: begin rgb_reg = 3'b011; end
            18'b001001001011011000: begin rgb_reg = 3'b001; end
            18'b001001001011011001: begin rgb_reg = 3'b011; end
            18'b001001001011011010: begin rgb_reg = 3'b011; end
            18'b001001001011011011: begin rgb_reg = 3'b011; end
            18'b001001001011100000: begin rgb_reg = 3'b011; end
            18'b001001001011100001: begin rgb_reg = 3'b011; end
            18'b001001001011100010: begin rgb_reg = 3'b011; end
            18'b001001001011100011: begin rgb_reg = 3'b011; end
            18'b001001001011110110: begin rgb_reg = 3'b001; end
            18'b001001001011110111: begin rgb_reg = 3'b011; end
            18'b001001001011111000: begin rgb_reg = 3'b011; end
            18'b001001001011111001: begin rgb_reg = 3'b011; end
            18'b001001001011111010: begin rgb_reg = 3'b001; end
            18'b001001001100000101: begin rgb_reg = 3'b001; end
            18'b001001001100000110: begin rgb_reg = 3'b011; end
            18'b001001001100000111: begin rgb_reg = 3'b011; end
            18'b001001001100001000: begin rgb_reg = 3'b011; end
            18'b001001001100001101: begin rgb_reg = 3'b011; end
            18'b001001001100001110: begin rgb_reg = 3'b011; end
            18'b001001001100001111: begin rgb_reg = 3'b011; end
            18'b001001001100010000: begin rgb_reg = 3'b011; end
            18'b001001001100011100: begin rgb_reg = 3'b011; end
            18'b001001001100011101: begin rgb_reg = 3'b011; end
            18'b001001001100011110: begin rgb_reg = 3'b011; end
            18'b001001001100011111: begin rgb_reg = 3'b011; end
            18'b001001001100100011: begin rgb_reg = 3'b001; end
            18'b001001001100100100: begin rgb_reg = 3'b011; end
            18'b001001001100100101: begin rgb_reg = 3'b011; end
            18'b001001001100100110: begin rgb_reg = 3'b011; end
            18'b001001001100100111: begin rgb_reg = 3'b001; end
            18'b001001001100110010: begin rgb_reg = 3'b001; end
            18'b001001001100110011: begin rgb_reg = 3'b011; end
            18'b001001001100110100: begin rgb_reg = 3'b011; end
            18'b001001001100110101: begin rgb_reg = 3'b011; end
            18'b001001001100111010: begin rgb_reg = 3'b011; end
            18'b001001001100111011: begin rgb_reg = 3'b011; end
            18'b001001001100111100: begin rgb_reg = 3'b011; end
            18'b001001001100111101: begin rgb_reg = 3'b011; end
            18'b001001001101001001: begin rgb_reg = 3'b011; end
            18'b001001001101001010: begin rgb_reg = 3'b011; end
            18'b001001001101001011: begin rgb_reg = 3'b011; end
            18'b001001001101001100: begin rgb_reg = 3'b001; end
            18'b001001001101010000: begin rgb_reg = 3'b001; end
            18'b001001001101010001: begin rgb_reg = 3'b011; end
            18'b001001001101010010: begin rgb_reg = 3'b011; end
            18'b001001001101010011: begin rgb_reg = 3'b011; end
            18'b001001001101010100: begin rgb_reg = 3'b001; end
            18'b001001010010011100: begin rgb_reg = 3'b001; end
            18'b001001010010011101: begin rgb_reg = 3'b011; end
            18'b001001010010011110: begin rgb_reg = 3'b011; end
            18'b001001010010011111: begin rgb_reg = 3'b011; end
            18'b001001010010101011: begin rgb_reg = 3'b001; end
            18'b001001010010101100: begin rgb_reg = 3'b011; end
            18'b001001010010101101: begin rgb_reg = 3'b011; end
            18'b001001010010101110: begin rgb_reg = 3'b011; end
            18'b001001010010110011: begin rgb_reg = 3'b011; end
            18'b001001010010110100: begin rgb_reg = 3'b011; end
            18'b001001010010110101: begin rgb_reg = 3'b011; end
            18'b001001010010110110: begin rgb_reg = 3'b011; end
            18'b001001010010111110: begin rgb_reg = 3'b011; end
            18'b001001010010111111: begin rgb_reg = 3'b011; end
            18'b001001010011000000: begin rgb_reg = 3'b011; end
            18'b001001010011000001: begin rgb_reg = 3'b011; end
            18'b001001010011000010: begin rgb_reg = 3'b011; end
            18'b001001010011000011: begin rgb_reg = 3'b011; end
            18'b001001010011000100: begin rgb_reg = 3'b011; end
            18'b001001010011000101: begin rgb_reg = 3'b011; end
            18'b001001010011001001: begin rgb_reg = 3'b001; end
            18'b001001010011001010: begin rgb_reg = 3'b011; end
            18'b001001010011001011: begin rgb_reg = 3'b011; end
            18'b001001010011001100: begin rgb_reg = 3'b011; end
            18'b001001010011011000: begin rgb_reg = 3'b001; end
            18'b001001010011011001: begin rgb_reg = 3'b011; end
            18'b001001010011011010: begin rgb_reg = 3'b011; end
            18'b001001010011011011: begin rgb_reg = 3'b011; end
            18'b001001010011100000: begin rgb_reg = 3'b011; end
            18'b001001010011100001: begin rgb_reg = 3'b011; end
            18'b001001010011100010: begin rgb_reg = 3'b011; end
            18'b001001010011100011: begin rgb_reg = 3'b011; end
            18'b001001010011110110: begin rgb_reg = 3'b001; end
            18'b001001010011110111: begin rgb_reg = 3'b011; end
            18'b001001010011111000: begin rgb_reg = 3'b011; end
            18'b001001010011111001: begin rgb_reg = 3'b011; end
            18'b001001010100000101: begin rgb_reg = 3'b001; end
            18'b001001010100000110: begin rgb_reg = 3'b011; end
            18'b001001010100000111: begin rgb_reg = 3'b011; end
            18'b001001010100001000: begin rgb_reg = 3'b011; end
            18'b001001010100001101: begin rgb_reg = 3'b011; end
            18'b001001010100001110: begin rgb_reg = 3'b011; end
            18'b001001010100001111: begin rgb_reg = 3'b011; end
            18'b001001010100010000: begin rgb_reg = 3'b011; end
            18'b001001010100011100: begin rgb_reg = 3'b011; end
            18'b001001010100011101: begin rgb_reg = 3'b011; end
            18'b001001010100011110: begin rgb_reg = 3'b011; end
            18'b001001010100011111: begin rgb_reg = 3'b011; end
            18'b001001010100100011: begin rgb_reg = 3'b001; end
            18'b001001010100100100: begin rgb_reg = 3'b011; end
            18'b001001010100100101: begin rgb_reg = 3'b011; end
            18'b001001010100100110: begin rgb_reg = 3'b011; end
            18'b001001010100110010: begin rgb_reg = 3'b001; end
            18'b001001010100110011: begin rgb_reg = 3'b011; end
            18'b001001010100110100: begin rgb_reg = 3'b011; end
            18'b001001010100110101: begin rgb_reg = 3'b011; end
            18'b001001010100111010: begin rgb_reg = 3'b011; end
            18'b001001010100111011: begin rgb_reg = 3'b011; end
            18'b001001010100111100: begin rgb_reg = 3'b011; end
            18'b001001010100111101: begin rgb_reg = 3'b011; end
            18'b001001010101001001: begin rgb_reg = 3'b011; end
            18'b001001010101001010: begin rgb_reg = 3'b011; end
            18'b001001010101001011: begin rgb_reg = 3'b011; end
            18'b001001010101001100: begin rgb_reg = 3'b011; end
            18'b001001010101010000: begin rgb_reg = 3'b001; end
            18'b001001010101010001: begin rgb_reg = 3'b011; end
            18'b001001010101010010: begin rgb_reg = 3'b011; end
            18'b001001010101010011: begin rgb_reg = 3'b011; end
            18'b001001011010011100: begin rgb_reg = 3'b001; end
            18'b001001011010011101: begin rgb_reg = 3'b011; end
            18'b001001011010011110: begin rgb_reg = 3'b011; end
            18'b001001011010011111: begin rgb_reg = 3'b011; end
            18'b001001011010101011: begin rgb_reg = 3'b001; end
            18'b001001011010101100: begin rgb_reg = 3'b011; end
            18'b001001011010101101: begin rgb_reg = 3'b011; end
            18'b001001011010101110: begin rgb_reg = 3'b011; end
            18'b001001011010110011: begin rgb_reg = 3'b011; end
            18'b001001011010110100: begin rgb_reg = 3'b011; end
            18'b001001011010110101: begin rgb_reg = 3'b011; end
            18'b001001011010110110: begin rgb_reg = 3'b011; end
            18'b001001011010111110: begin rgb_reg = 3'b011; end
            18'b001001011010111111: begin rgb_reg = 3'b011; end
            18'b001001011011000000: begin rgb_reg = 3'b011; end
            18'b001001011011000001: begin rgb_reg = 3'b011; end
            18'b001001011011000010: begin rgb_reg = 3'b011; end
            18'b001001011011000011: begin rgb_reg = 3'b011; end
            18'b001001011011000100: begin rgb_reg = 3'b011; end
            18'b001001011011000101: begin rgb_reg = 3'b011; end
            18'b001001011011001001: begin rgb_reg = 3'b001; end
            18'b001001011011001010: begin rgb_reg = 3'b011; end
            18'b001001011011001011: begin rgb_reg = 3'b011; end
            18'b001001011011001100: begin rgb_reg = 3'b011; end
            18'b001001011011011000: begin rgb_reg = 3'b001; end
            18'b001001011011011001: begin rgb_reg = 3'b011; end
            18'b001001011011011010: begin rgb_reg = 3'b011; end
            18'b001001011011011011: begin rgb_reg = 3'b011; end
            18'b001001011011100000: begin rgb_reg = 3'b011; end
            18'b001001011011100001: begin rgb_reg = 3'b011; end
            18'b001001011011100010: begin rgb_reg = 3'b011; end
            18'b001001011011100011: begin rgb_reg = 3'b011; end
            18'b001001011011110110: begin rgb_reg = 3'b001; end
            18'b001001011011110111: begin rgb_reg = 3'b011; end
            18'b001001011011111000: begin rgb_reg = 3'b011; end
            18'b001001011011111001: begin rgb_reg = 3'b011; end
            18'b001001011100000101: begin rgb_reg = 3'b001; end
            18'b001001011100000110: begin rgb_reg = 3'b011; end
            18'b001001011100000111: begin rgb_reg = 3'b011; end
            18'b001001011100001000: begin rgb_reg = 3'b011; end
            18'b001001011100001101: begin rgb_reg = 3'b011; end
            18'b001001011100001110: begin rgb_reg = 3'b011; end
            18'b001001011100001111: begin rgb_reg = 3'b011; end
            18'b001001011100010000: begin rgb_reg = 3'b011; end
            18'b001001011100011100: begin rgb_reg = 3'b011; end
            18'b001001011100011101: begin rgb_reg = 3'b011; end
            18'b001001011100011110: begin rgb_reg = 3'b011; end
            18'b001001011100011111: begin rgb_reg = 3'b011; end
            18'b001001011100100011: begin rgb_reg = 3'b001; end
            18'b001001011100100100: begin rgb_reg = 3'b011; end
            18'b001001011100100101: begin rgb_reg = 3'b011; end
            18'b001001011100100110: begin rgb_reg = 3'b011; end
            18'b001001011100110010: begin rgb_reg = 3'b001; end
            18'b001001011100110011: begin rgb_reg = 3'b011; end
            18'b001001011100110100: begin rgb_reg = 3'b011; end
            18'b001001011100110101: begin rgb_reg = 3'b011; end
            18'b001001011100111010: begin rgb_reg = 3'b011; end
            18'b001001011100111011: begin rgb_reg = 3'b011; end
            18'b001001011100111100: begin rgb_reg = 3'b011; end
            18'b001001011100111101: begin rgb_reg = 3'b011; end
            18'b001001011101001001: begin rgb_reg = 3'b011; end
            18'b001001011101001010: begin rgb_reg = 3'b011; end
            18'b001001011101001011: begin rgb_reg = 3'b011; end
            18'b001001011101001100: begin rgb_reg = 3'b011; end
            18'b001001011101010000: begin rgb_reg = 3'b001; end
            18'b001001011101010001: begin rgb_reg = 3'b011; end
            18'b001001011101010010: begin rgb_reg = 3'b011; end
            18'b001001011101010011: begin rgb_reg = 3'b011; end
            18'b001001100010011100: begin rgb_reg = 3'b001; end
            18'b001001100010011101: begin rgb_reg = 3'b011; end
            18'b001001100010011110: begin rgb_reg = 3'b011; end
            18'b001001100010011111: begin rgb_reg = 3'b011; end
            18'b001001100010101011: begin rgb_reg = 3'b001; end
            18'b001001100010101100: begin rgb_reg = 3'b011; end
            18'b001001100010101101: begin rgb_reg = 3'b011; end
            18'b001001100010101110: begin rgb_reg = 3'b011; end
            18'b001001100010110011: begin rgb_reg = 3'b011; end
            18'b001001100010110100: begin rgb_reg = 3'b011; end
            18'b001001100010110101: begin rgb_reg = 3'b011; end
            18'b001001100010110110: begin rgb_reg = 3'b011; end
            18'b001001100010111110: begin rgb_reg = 3'b011; end
            18'b001001100010111111: begin rgb_reg = 3'b011; end
            18'b001001100011000000: begin rgb_reg = 3'b011; end
            18'b001001100011000001: begin rgb_reg = 3'b011; end
            18'b001001100011000010: begin rgb_reg = 3'b011; end
            18'b001001100011000011: begin rgb_reg = 3'b011; end
            18'b001001100011000100: begin rgb_reg = 3'b011; end
            18'b001001100011000101: begin rgb_reg = 3'b011; end
            18'b001001100011001001: begin rgb_reg = 3'b001; end
            18'b001001100011001010: begin rgb_reg = 3'b011; end
            18'b001001100011001011: begin rgb_reg = 3'b011; end
            18'b001001100011001100: begin rgb_reg = 3'b011; end
            18'b001001100011011000: begin rgb_reg = 3'b001; end
            18'b001001100011011001: begin rgb_reg = 3'b011; end
            18'b001001100011011010: begin rgb_reg = 3'b011; end
            18'b001001100011011011: begin rgb_reg = 3'b011; end
            18'b001001100011100000: begin rgb_reg = 3'b011; end
            18'b001001100011100001: begin rgb_reg = 3'b011; end
            18'b001001100011100010: begin rgb_reg = 3'b011; end
            18'b001001100011100011: begin rgb_reg = 3'b011; end
            18'b001001100011110110: begin rgb_reg = 3'b001; end
            18'b001001100011110111: begin rgb_reg = 3'b011; end
            18'b001001100011111000: begin rgb_reg = 3'b011; end
            18'b001001100011111001: begin rgb_reg = 3'b011; end
            18'b001001100100000101: begin rgb_reg = 3'b001; end
            18'b001001100100000110: begin rgb_reg = 3'b011; end
            18'b001001100100000111: begin rgb_reg = 3'b011; end
            18'b001001100100001000: begin rgb_reg = 3'b011; end
            18'b001001100100001101: begin rgb_reg = 3'b011; end
            18'b001001100100001110: begin rgb_reg = 3'b011; end
            18'b001001100100001111: begin rgb_reg = 3'b011; end
            18'b001001100100010000: begin rgb_reg = 3'b011; end
            18'b001001100100011100: begin rgb_reg = 3'b011; end
            18'b001001100100011101: begin rgb_reg = 3'b011; end
            18'b001001100100011110: begin rgb_reg = 3'b011; end
            18'b001001100100011111: begin rgb_reg = 3'b011; end
            18'b001001100100100011: begin rgb_reg = 3'b001; end
            18'b001001100100100100: begin rgb_reg = 3'b011; end
            18'b001001100100100101: begin rgb_reg = 3'b011; end
            18'b001001100100100110: begin rgb_reg = 3'b011; end
            18'b001001100100110010: begin rgb_reg = 3'b001; end
            18'b001001100100110011: begin rgb_reg = 3'b011; end
            18'b001001100100110100: begin rgb_reg = 3'b011; end
            18'b001001100100110101: begin rgb_reg = 3'b011; end
            18'b001001100100111010: begin rgb_reg = 3'b011; end
            18'b001001100100111011: begin rgb_reg = 3'b011; end
            18'b001001100100111100: begin rgb_reg = 3'b011; end
            18'b001001100100111101: begin rgb_reg = 3'b011; end
            18'b001001100101001001: begin rgb_reg = 3'b011; end
            18'b001001100101001010: begin rgb_reg = 3'b011; end
            18'b001001100101001011: begin rgb_reg = 3'b011; end
            18'b001001100101001100: begin rgb_reg = 3'b011; end
            18'b001001100101010000: begin rgb_reg = 3'b001; end
            18'b001001100101010001: begin rgb_reg = 3'b011; end
            18'b001001100101010010: begin rgb_reg = 3'b011; end
            18'b001001100101010011: begin rgb_reg = 3'b011; end
            18'b001001101010011100: begin rgb_reg = 3'b001; end
            18'b001001101010011101: begin rgb_reg = 3'b011; end
            18'b001001101010011110: begin rgb_reg = 3'b011; end
            18'b001001101010011111: begin rgb_reg = 3'b011; end
            18'b001001101010101011: begin rgb_reg = 3'b001; end
            18'b001001101010101100: begin rgb_reg = 3'b011; end
            18'b001001101010101101: begin rgb_reg = 3'b011; end
            18'b001001101010101110: begin rgb_reg = 3'b011; end
            18'b001001101010110011: begin rgb_reg = 3'b011; end
            18'b001001101010110100: begin rgb_reg = 3'b011; end
            18'b001001101010110101: begin rgb_reg = 3'b011; end
            18'b001001101010110110: begin rgb_reg = 3'b011; end
            18'b001001101011000010: begin rgb_reg = 3'b011; end
            18'b001001101011000011: begin rgb_reg = 3'b011; end
            18'b001001101011000100: begin rgb_reg = 3'b011; end
            18'b001001101011000101: begin rgb_reg = 3'b011; end
            18'b001001101011001001: begin rgb_reg = 3'b001; end
            18'b001001101011001010: begin rgb_reg = 3'b011; end
            18'b001001101011001011: begin rgb_reg = 3'b011; end
            18'b001001101011001100: begin rgb_reg = 3'b011; end
            18'b001001101011011000: begin rgb_reg = 3'b001; end
            18'b001001101011011001: begin rgb_reg = 3'b011; end
            18'b001001101011011010: begin rgb_reg = 3'b011; end
            18'b001001101011011011: begin rgb_reg = 3'b011; end
            18'b001001101011100000: begin rgb_reg = 3'b011; end
            18'b001001101011100001: begin rgb_reg = 3'b011; end
            18'b001001101011100010: begin rgb_reg = 3'b011; end
            18'b001001101011100011: begin rgb_reg = 3'b011; end
            18'b001001101011110110: begin rgb_reg = 3'b001; end
            18'b001001101011110111: begin rgb_reg = 3'b011; end
            18'b001001101011111000: begin rgb_reg = 3'b011; end
            18'b001001101011111001: begin rgb_reg = 3'b011; end
            18'b001001101100000101: begin rgb_reg = 3'b001; end
            18'b001001101100000110: begin rgb_reg = 3'b011; end
            18'b001001101100000111: begin rgb_reg = 3'b011; end
            18'b001001101100001000: begin rgb_reg = 3'b011; end
            18'b001001101100001101: begin rgb_reg = 3'b011; end
            18'b001001101100001110: begin rgb_reg = 3'b011; end
            18'b001001101100001111: begin rgb_reg = 3'b011; end
            18'b001001101100010000: begin rgb_reg = 3'b011; end
            18'b001001101100010100: begin rgb_reg = 3'b001; end
            18'b001001101100010101: begin rgb_reg = 3'b011; end
            18'b001001101100010110: begin rgb_reg = 3'b011; end
            18'b001001101100010111: begin rgb_reg = 3'b011; end
            18'b001001101100011100: begin rgb_reg = 3'b011; end
            18'b001001101100011101: begin rgb_reg = 3'b011; end
            18'b001001101100011110: begin rgb_reg = 3'b011; end
            18'b001001101100011111: begin rgb_reg = 3'b011; end
            18'b001001101100100011: begin rgb_reg = 3'b001; end
            18'b001001101100100100: begin rgb_reg = 3'b011; end
            18'b001001101100100101: begin rgb_reg = 3'b011; end
            18'b001001101100100110: begin rgb_reg = 3'b011; end
            18'b001001101100110010: begin rgb_reg = 3'b001; end
            18'b001001101100110011: begin rgb_reg = 3'b011; end
            18'b001001101100110100: begin rgb_reg = 3'b011; end
            18'b001001101100110101: begin rgb_reg = 3'b011; end
            18'b001001101100111010: begin rgb_reg = 3'b011; end
            18'b001001101100111011: begin rgb_reg = 3'b011; end
            18'b001001101100111100: begin rgb_reg = 3'b011; end
            18'b001001101100111101: begin rgb_reg = 3'b011; end
            18'b001001101101001001: begin rgb_reg = 3'b011; end
            18'b001001101101001010: begin rgb_reg = 3'b011; end
            18'b001001101101001011: begin rgb_reg = 3'b011; end
            18'b001001101101001100: begin rgb_reg = 3'b011; end
            18'b001001101101010000: begin rgb_reg = 3'b001; end
            18'b001001101101010001: begin rgb_reg = 3'b011; end
            18'b001001101101010010: begin rgb_reg = 3'b011; end
            18'b001001101101010011: begin rgb_reg = 3'b011; end
            18'b001001110010011100: begin rgb_reg = 3'b001; end
            18'b001001110010011101: begin rgb_reg = 3'b011; end
            18'b001001110010011110: begin rgb_reg = 3'b011; end
            18'b001001110010011111: begin rgb_reg = 3'b011; end
            18'b001001110010101011: begin rgb_reg = 3'b001; end
            18'b001001110010101100: begin rgb_reg = 3'b011; end
            18'b001001110010101101: begin rgb_reg = 3'b011; end
            18'b001001110010101110: begin rgb_reg = 3'b011; end
            18'b001001110010110011: begin rgb_reg = 3'b011; end
            18'b001001110010110100: begin rgb_reg = 3'b011; end
            18'b001001110010110101: begin rgb_reg = 3'b011; end
            18'b001001110010110110: begin rgb_reg = 3'b011; end
            18'b001001110011000010: begin rgb_reg = 3'b011; end
            18'b001001110011000011: begin rgb_reg = 3'b011; end
            18'b001001110011000100: begin rgb_reg = 3'b011; end
            18'b001001110011000101: begin rgb_reg = 3'b011; end
            18'b001001110011001001: begin rgb_reg = 3'b001; end
            18'b001001110011001010: begin rgb_reg = 3'b011; end
            18'b001001110011001011: begin rgb_reg = 3'b011; end
            18'b001001110011001100: begin rgb_reg = 3'b011; end
            18'b001001110011011000: begin rgb_reg = 3'b001; end
            18'b001001110011011001: begin rgb_reg = 3'b011; end
            18'b001001110011011010: begin rgb_reg = 3'b011; end
            18'b001001110011011011: begin rgb_reg = 3'b011; end
            18'b001001110011100000: begin rgb_reg = 3'b011; end
            18'b001001110011100001: begin rgb_reg = 3'b011; end
            18'b001001110011100010: begin rgb_reg = 3'b011; end
            18'b001001110011100011: begin rgb_reg = 3'b011; end
            18'b001001110011110110: begin rgb_reg = 3'b001; end
            18'b001001110011110111: begin rgb_reg = 3'b011; end
            18'b001001110011111000: begin rgb_reg = 3'b011; end
            18'b001001110011111001: begin rgb_reg = 3'b011; end
            18'b001001110100000101: begin rgb_reg = 3'b001; end
            18'b001001110100000110: begin rgb_reg = 3'b011; end
            18'b001001110100000111: begin rgb_reg = 3'b011; end
            18'b001001110100001000: begin rgb_reg = 3'b011; end
            18'b001001110100001101: begin rgb_reg = 3'b011; end
            18'b001001110100001110: begin rgb_reg = 3'b011; end
            18'b001001110100001111: begin rgb_reg = 3'b011; end
            18'b001001110100010000: begin rgb_reg = 3'b011; end
            18'b001001110100010100: begin rgb_reg = 3'b001; end
            18'b001001110100010101: begin rgb_reg = 3'b011; end
            18'b001001110100010110: begin rgb_reg = 3'b011; end
            18'b001001110100010111: begin rgb_reg = 3'b011; end
            18'b001001110100011100: begin rgb_reg = 3'b011; end
            18'b001001110100011101: begin rgb_reg = 3'b011; end
            18'b001001110100011110: begin rgb_reg = 3'b011; end
            18'b001001110100011111: begin rgb_reg = 3'b011; end
            18'b001001110100100011: begin rgb_reg = 3'b001; end
            18'b001001110100100100: begin rgb_reg = 3'b011; end
            18'b001001110100100101: begin rgb_reg = 3'b011; end
            18'b001001110100100110: begin rgb_reg = 3'b011; end
            18'b001001110100110010: begin rgb_reg = 3'b001; end
            18'b001001110100110011: begin rgb_reg = 3'b011; end
            18'b001001110100110100: begin rgb_reg = 3'b011; end
            18'b001001110100110101: begin rgb_reg = 3'b011; end
            18'b001001110100111010: begin rgb_reg = 3'b011; end
            18'b001001110100111011: begin rgb_reg = 3'b011; end
            18'b001001110100111100: begin rgb_reg = 3'b011; end
            18'b001001110100111101: begin rgb_reg = 3'b011; end
            18'b001001110101001001: begin rgb_reg = 3'b011; end
            18'b001001110101001010: begin rgb_reg = 3'b011; end
            18'b001001110101001011: begin rgb_reg = 3'b011; end
            18'b001001110101001100: begin rgb_reg = 3'b011; end
            18'b001001110101010000: begin rgb_reg = 3'b001; end
            18'b001001110101010001: begin rgb_reg = 3'b011; end
            18'b001001110101010010: begin rgb_reg = 3'b011; end
            18'b001001110101010011: begin rgb_reg = 3'b011; end
            18'b001001111010011100: begin rgb_reg = 3'b001; end
            18'b001001111010011101: begin rgb_reg = 3'b011; end
            18'b001001111010011110: begin rgb_reg = 3'b011; end
            18'b001001111010011111: begin rgb_reg = 3'b011; end
            18'b001001111010101011: begin rgb_reg = 3'b001; end
            18'b001001111010101100: begin rgb_reg = 3'b011; end
            18'b001001111010101101: begin rgb_reg = 3'b011; end
            18'b001001111010101110: begin rgb_reg = 3'b011; end
            18'b001001111010110011: begin rgb_reg = 3'b011; end
            18'b001001111010110100: begin rgb_reg = 3'b011; end
            18'b001001111010110101: begin rgb_reg = 3'b011; end
            18'b001001111010110110: begin rgb_reg = 3'b011; end
            18'b001001111011000010: begin rgb_reg = 3'b011; end
            18'b001001111011000011: begin rgb_reg = 3'b011; end
            18'b001001111011000100: begin rgb_reg = 3'b011; end
            18'b001001111011000101: begin rgb_reg = 3'b011; end
            18'b001001111011001001: begin rgb_reg = 3'b001; end
            18'b001001111011001010: begin rgb_reg = 3'b011; end
            18'b001001111011001011: begin rgb_reg = 3'b011; end
            18'b001001111011001100: begin rgb_reg = 3'b011; end
            18'b001001111011011000: begin rgb_reg = 3'b001; end
            18'b001001111011011001: begin rgb_reg = 3'b011; end
            18'b001001111011011010: begin rgb_reg = 3'b011; end
            18'b001001111011011011: begin rgb_reg = 3'b011; end
            18'b001001111011100000: begin rgb_reg = 3'b011; end
            18'b001001111011100001: begin rgb_reg = 3'b011; end
            18'b001001111011100010: begin rgb_reg = 3'b011; end
            18'b001001111011100011: begin rgb_reg = 3'b011; end
            18'b001001111011110110: begin rgb_reg = 3'b001; end
            18'b001001111011110111: begin rgb_reg = 3'b011; end
            18'b001001111011111000: begin rgb_reg = 3'b011; end
            18'b001001111011111001: begin rgb_reg = 3'b011; end
            18'b001001111100000101: begin rgb_reg = 3'b001; end
            18'b001001111100000110: begin rgb_reg = 3'b011; end
            18'b001001111100000111: begin rgb_reg = 3'b011; end
            18'b001001111100001000: begin rgb_reg = 3'b011; end
            18'b001001111100001101: begin rgb_reg = 3'b011; end
            18'b001001111100001110: begin rgb_reg = 3'b011; end
            18'b001001111100001111: begin rgb_reg = 3'b011; end
            18'b001001111100010000: begin rgb_reg = 3'b011; end
            18'b001001111100010100: begin rgb_reg = 3'b001; end
            18'b001001111100010101: begin rgb_reg = 3'b011; end
            18'b001001111100010110: begin rgb_reg = 3'b011; end
            18'b001001111100010111: begin rgb_reg = 3'b011; end
            18'b001001111100011100: begin rgb_reg = 3'b011; end
            18'b001001111100011101: begin rgb_reg = 3'b011; end
            18'b001001111100011110: begin rgb_reg = 3'b011; end
            18'b001001111100011111: begin rgb_reg = 3'b011; end
            18'b001001111100100011: begin rgb_reg = 3'b001; end
            18'b001001111100100100: begin rgb_reg = 3'b011; end
            18'b001001111100100101: begin rgb_reg = 3'b011; end
            18'b001001111100100110: begin rgb_reg = 3'b011; end
            18'b001001111100110010: begin rgb_reg = 3'b001; end
            18'b001001111100110011: begin rgb_reg = 3'b011; end
            18'b001001111100110100: begin rgb_reg = 3'b011; end
            18'b001001111100110101: begin rgb_reg = 3'b011; end
            18'b001001111100111010: begin rgb_reg = 3'b011; end
            18'b001001111100111011: begin rgb_reg = 3'b011; end
            18'b001001111100111100: begin rgb_reg = 3'b011; end
            18'b001001111100111101: begin rgb_reg = 3'b011; end
            18'b001001111101001001: begin rgb_reg = 3'b011; end
            18'b001001111101001010: begin rgb_reg = 3'b011; end
            18'b001001111101001011: begin rgb_reg = 3'b011; end
            18'b001001111101001100: begin rgb_reg = 3'b011; end
            18'b001001111101010000: begin rgb_reg = 3'b001; end
            18'b001001111101010001: begin rgb_reg = 3'b011; end
            18'b001001111101010010: begin rgb_reg = 3'b011; end
            18'b001001111101010011: begin rgb_reg = 3'b011; end
            18'b001010000010011100: begin rgb_reg = 3'b001; end
            18'b001010000010011101: begin rgb_reg = 3'b011; end
            18'b001010000010011110: begin rgb_reg = 3'b011; end
            18'b001010000010011111: begin rgb_reg = 3'b011; end
            18'b001010000010101011: begin rgb_reg = 3'b001; end
            18'b001010000010101100: begin rgb_reg = 3'b011; end
            18'b001010000010101101: begin rgb_reg = 3'b011; end
            18'b001010000010101110: begin rgb_reg = 3'b011; end
            18'b001010000010110011: begin rgb_reg = 3'b011; end
            18'b001010000010110100: begin rgb_reg = 3'b011; end
            18'b001010000010110101: begin rgb_reg = 3'b011; end
            18'b001010000010110110: begin rgb_reg = 3'b011; end
            18'b001010000011000010: begin rgb_reg = 3'b011; end
            18'b001010000011000011: begin rgb_reg = 3'b011; end
            18'b001010000011000100: begin rgb_reg = 3'b011; end
            18'b001010000011000101: begin rgb_reg = 3'b011; end
            18'b001010000011001001: begin rgb_reg = 3'b001; end
            18'b001010000011001010: begin rgb_reg = 3'b011; end
            18'b001010000011001011: begin rgb_reg = 3'b011; end
            18'b001010000011001100: begin rgb_reg = 3'b011; end
            18'b001010000011011000: begin rgb_reg = 3'b001; end
            18'b001010000011011001: begin rgb_reg = 3'b011; end
            18'b001010000011011010: begin rgb_reg = 3'b011; end
            18'b001010000011011011: begin rgb_reg = 3'b011; end
            18'b001010000011100000: begin rgb_reg = 3'b011; end
            18'b001010000011100001: begin rgb_reg = 3'b011; end
            18'b001010000011100010: begin rgb_reg = 3'b011; end
            18'b001010000011100011: begin rgb_reg = 3'b011; end
            18'b001010000011110110: begin rgb_reg = 3'b001; end
            18'b001010000011110111: begin rgb_reg = 3'b011; end
            18'b001010000011111000: begin rgb_reg = 3'b011; end
            18'b001010000011111001: begin rgb_reg = 3'b011; end
            18'b001010000100000101: begin rgb_reg = 3'b001; end
            18'b001010000100000110: begin rgb_reg = 3'b011; end
            18'b001010000100000111: begin rgb_reg = 3'b011; end
            18'b001010000100001000: begin rgb_reg = 3'b011; end
            18'b001010000100001101: begin rgb_reg = 3'b011; end
            18'b001010000100001110: begin rgb_reg = 3'b011; end
            18'b001010000100001111: begin rgb_reg = 3'b011; end
            18'b001010000100010000: begin rgb_reg = 3'b011; end
            18'b001010000100010100: begin rgb_reg = 3'b001; end
            18'b001010000100010101: begin rgb_reg = 3'b011; end
            18'b001010000100010110: begin rgb_reg = 3'b011; end
            18'b001010000100010111: begin rgb_reg = 3'b011; end
            18'b001010000100011000: begin rgb_reg = 3'b001; end
            18'b001010000100011100: begin rgb_reg = 3'b011; end
            18'b001010000100011101: begin rgb_reg = 3'b011; end
            18'b001010000100011110: begin rgb_reg = 3'b011; end
            18'b001010000100011111: begin rgb_reg = 3'b011; end
            18'b001010000100100011: begin rgb_reg = 3'b001; end
            18'b001010000100100100: begin rgb_reg = 3'b011; end
            18'b001010000100100101: begin rgb_reg = 3'b011; end
            18'b001010000100100110: begin rgb_reg = 3'b011; end
            18'b001010000100110010: begin rgb_reg = 3'b001; end
            18'b001010000100110011: begin rgb_reg = 3'b011; end
            18'b001010000100110100: begin rgb_reg = 3'b011; end
            18'b001010000100110101: begin rgb_reg = 3'b011; end
            18'b001010000100111010: begin rgb_reg = 3'b011; end
            18'b001010000100111011: begin rgb_reg = 3'b011; end
            18'b001010000100111100: begin rgb_reg = 3'b011; end
            18'b001010000100111101: begin rgb_reg = 3'b011; end
            18'b001010000101001001: begin rgb_reg = 3'b011; end
            18'b001010000101001010: begin rgb_reg = 3'b011; end
            18'b001010000101001011: begin rgb_reg = 3'b011; end
            18'b001010000101001100: begin rgb_reg = 3'b011; end
            18'b001010000101010000: begin rgb_reg = 3'b001; end
            18'b001010000101010001: begin rgb_reg = 3'b011; end
            18'b001010000101010010: begin rgb_reg = 3'b011; end
            18'b001010000101010011: begin rgb_reg = 3'b011; end
            18'b001010001010011100: begin rgb_reg = 3'b001; end
            18'b001010001010011101: begin rgb_reg = 3'b011; end
            18'b001010001010011110: begin rgb_reg = 3'b011; end
            18'b001010001010011111: begin rgb_reg = 3'b011; end
            18'b001010001010101011: begin rgb_reg = 3'b001; end
            18'b001010001010101100: begin rgb_reg = 3'b011; end
            18'b001010001010101101: begin rgb_reg = 3'b011; end
            18'b001010001010101110: begin rgb_reg = 3'b011; end
            18'b001010001010110011: begin rgb_reg = 3'b011; end
            18'b001010001010110100: begin rgb_reg = 3'b011; end
            18'b001010001010110101: begin rgb_reg = 3'b011; end
            18'b001010001010110110: begin rgb_reg = 3'b011; end
            18'b001010001011000010: begin rgb_reg = 3'b011; end
            18'b001010001011000011: begin rgb_reg = 3'b011; end
            18'b001010001011000100: begin rgb_reg = 3'b011; end
            18'b001010001011000101: begin rgb_reg = 3'b011; end
            18'b001010001011001001: begin rgb_reg = 3'b001; end
            18'b001010001011001010: begin rgb_reg = 3'b011; end
            18'b001010001011001011: begin rgb_reg = 3'b011; end
            18'b001010001011001100: begin rgb_reg = 3'b011; end
            18'b001010001011011000: begin rgb_reg = 3'b001; end
            18'b001010001011011001: begin rgb_reg = 3'b011; end
            18'b001010001011011010: begin rgb_reg = 3'b011; end
            18'b001010001011011011: begin rgb_reg = 3'b011; end
            18'b001010001011100000: begin rgb_reg = 3'b011; end
            18'b001010001011100001: begin rgb_reg = 3'b011; end
            18'b001010001011100010: begin rgb_reg = 3'b011; end
            18'b001010001011100011: begin rgb_reg = 3'b011; end
            18'b001010001011110110: begin rgb_reg = 3'b001; end
            18'b001010001011110111: begin rgb_reg = 3'b011; end
            18'b001010001011111000: begin rgb_reg = 3'b011; end
            18'b001010001011111001: begin rgb_reg = 3'b011; end
            18'b001010001100000101: begin rgb_reg = 3'b001; end
            18'b001010001100000110: begin rgb_reg = 3'b011; end
            18'b001010001100000111: begin rgb_reg = 3'b011; end
            18'b001010001100001000: begin rgb_reg = 3'b011; end
            18'b001010001100001101: begin rgb_reg = 3'b011; end
            18'b001010001100001110: begin rgb_reg = 3'b011; end
            18'b001010001100001111: begin rgb_reg = 3'b011; end
            18'b001010001100010000: begin rgb_reg = 3'b011; end
            18'b001010001100010001: begin rgb_reg = 3'b011; end
            18'b001010001100010010: begin rgb_reg = 3'b011; end
            18'b001010001100010011: begin rgb_reg = 3'b011; end
            18'b001010001100010100: begin rgb_reg = 3'b001; end
            18'b001010001100011000: begin rgb_reg = 3'b011; end
            18'b001010001100011001: begin rgb_reg = 3'b011; end
            18'b001010001100011010: begin rgb_reg = 3'b011; end
            18'b001010001100011011: begin rgb_reg = 3'b011; end
            18'b001010001100011100: begin rgb_reg = 3'b011; end
            18'b001010001100011101: begin rgb_reg = 3'b011; end
            18'b001010001100011110: begin rgb_reg = 3'b011; end
            18'b001010001100011111: begin rgb_reg = 3'b011; end
            18'b001010001100100011: begin rgb_reg = 3'b001; end
            18'b001010001100100100: begin rgb_reg = 3'b011; end
            18'b001010001100100101: begin rgb_reg = 3'b011; end
            18'b001010001100100110: begin rgb_reg = 3'b011; end
            18'b001010001100110010: begin rgb_reg = 3'b001; end
            18'b001010001100110011: begin rgb_reg = 3'b011; end
            18'b001010001100110100: begin rgb_reg = 3'b011; end
            18'b001010001100110101: begin rgb_reg = 3'b011; end
            18'b001010001100111010: begin rgb_reg = 3'b011; end
            18'b001010001100111011: begin rgb_reg = 3'b011; end
            18'b001010001100111100: begin rgb_reg = 3'b011; end
            18'b001010001100111101: begin rgb_reg = 3'b011; end
            18'b001010001101001001: begin rgb_reg = 3'b011; end
            18'b001010001101001010: begin rgb_reg = 3'b011; end
            18'b001010001101001011: begin rgb_reg = 3'b011; end
            18'b001010001101001100: begin rgb_reg = 3'b011; end
            18'b001010001101010000: begin rgb_reg = 3'b001; end
            18'b001010001101010001: begin rgb_reg = 3'b011; end
            18'b001010001101010010: begin rgb_reg = 3'b011; end
            18'b001010001101010011: begin rgb_reg = 3'b011; end
            18'b001010010010011100: begin rgb_reg = 3'b001; end
            18'b001010010010011101: begin rgb_reg = 3'b011; end
            18'b001010010010011110: begin rgb_reg = 3'b011; end
            18'b001010010010011111: begin rgb_reg = 3'b011; end
            18'b001010010010101011: begin rgb_reg = 3'b001; end
            18'b001010010010101100: begin rgb_reg = 3'b011; end
            18'b001010010010101101: begin rgb_reg = 3'b011; end
            18'b001010010010101110: begin rgb_reg = 3'b011; end
            18'b001010010010110011: begin rgb_reg = 3'b011; end
            18'b001010010010110100: begin rgb_reg = 3'b011; end
            18'b001010010010110101: begin rgb_reg = 3'b011; end
            18'b001010010010110110: begin rgb_reg = 3'b011; end
            18'b001010010011000010: begin rgb_reg = 3'b011; end
            18'b001010010011000011: begin rgb_reg = 3'b011; end
            18'b001010010011000100: begin rgb_reg = 3'b011; end
            18'b001010010011000101: begin rgb_reg = 3'b011; end
            18'b001010010011001001: begin rgb_reg = 3'b001; end
            18'b001010010011001010: begin rgb_reg = 3'b011; end
            18'b001010010011001011: begin rgb_reg = 3'b011; end
            18'b001010010011001100: begin rgb_reg = 3'b011; end
            18'b001010010011011000: begin rgb_reg = 3'b001; end
            18'b001010010011011001: begin rgb_reg = 3'b011; end
            18'b001010010011011010: begin rgb_reg = 3'b011; end
            18'b001010010011011011: begin rgb_reg = 3'b011; end
            18'b001010010011100000: begin rgb_reg = 3'b011; end
            18'b001010010011100001: begin rgb_reg = 3'b011; end
            18'b001010010011100010: begin rgb_reg = 3'b011; end
            18'b001010010011100011: begin rgb_reg = 3'b011; end
            18'b001010010011110110: begin rgb_reg = 3'b001; end
            18'b001010010011110111: begin rgb_reg = 3'b011; end
            18'b001010010011111000: begin rgb_reg = 3'b011; end
            18'b001010010011111001: begin rgb_reg = 3'b011; end
            18'b001010010100000101: begin rgb_reg = 3'b001; end
            18'b001010010100000110: begin rgb_reg = 3'b011; end
            18'b001010010100000111: begin rgb_reg = 3'b011; end
            18'b001010010100001000: begin rgb_reg = 3'b011; end
            18'b001010010100001101: begin rgb_reg = 3'b011; end
            18'b001010010100001110: begin rgb_reg = 3'b011; end
            18'b001010010100001111: begin rgb_reg = 3'b011; end
            18'b001010010100010000: begin rgb_reg = 3'b011; end
            18'b001010010100010001: begin rgb_reg = 3'b011; end
            18'b001010010100010010: begin rgb_reg = 3'b011; end
            18'b001010010100010011: begin rgb_reg = 3'b011; end
            18'b001010010100010100: begin rgb_reg = 3'b001; end
            18'b001010010100011000: begin rgb_reg = 3'b011; end
            18'b001010010100011001: begin rgb_reg = 3'b011; end
            18'b001010010100011010: begin rgb_reg = 3'b011; end
            18'b001010010100011011: begin rgb_reg = 3'b011; end
            18'b001010010100011100: begin rgb_reg = 3'b011; end
            18'b001010010100011101: begin rgb_reg = 3'b011; end
            18'b001010010100011110: begin rgb_reg = 3'b011; end
            18'b001010010100011111: begin rgb_reg = 3'b011; end
            18'b001010010100100011: begin rgb_reg = 3'b001; end
            18'b001010010100100100: begin rgb_reg = 3'b011; end
            18'b001010010100100101: begin rgb_reg = 3'b011; end
            18'b001010010100100110: begin rgb_reg = 3'b011; end
            18'b001010010100110010: begin rgb_reg = 3'b001; end
            18'b001010010100110011: begin rgb_reg = 3'b011; end
            18'b001010010100110100: begin rgb_reg = 3'b011; end
            18'b001010010100110101: begin rgb_reg = 3'b011; end
            18'b001010010100111010: begin rgb_reg = 3'b011; end
            18'b001010010100111011: begin rgb_reg = 3'b011; end
            18'b001010010100111100: begin rgb_reg = 3'b011; end
            18'b001010010100111101: begin rgb_reg = 3'b011; end
            18'b001010010101001001: begin rgb_reg = 3'b011; end
            18'b001010010101001010: begin rgb_reg = 3'b011; end
            18'b001010010101001011: begin rgb_reg = 3'b011; end
            18'b001010010101001100: begin rgb_reg = 3'b011; end
            18'b001010010101010000: begin rgb_reg = 3'b001; end
            18'b001010010101010001: begin rgb_reg = 3'b011; end
            18'b001010010101010010: begin rgb_reg = 3'b011; end
            18'b001010010101010011: begin rgb_reg = 3'b011; end
            18'b001010011010011100: begin rgb_reg = 3'b001; end
            18'b001010011010011101: begin rgb_reg = 3'b011; end
            18'b001010011010011110: begin rgb_reg = 3'b011; end
            18'b001010011010011111: begin rgb_reg = 3'b011; end
            18'b001010011010101011: begin rgb_reg = 3'b001; end
            18'b001010011010101100: begin rgb_reg = 3'b011; end
            18'b001010011010101101: begin rgb_reg = 3'b011; end
            18'b001010011010101110: begin rgb_reg = 3'b011; end
            18'b001010011010110011: begin rgb_reg = 3'b011; end
            18'b001010011010110100: begin rgb_reg = 3'b011; end
            18'b001010011010110101: begin rgb_reg = 3'b011; end
            18'b001010011010110110: begin rgb_reg = 3'b011; end
            18'b001010011011000010: begin rgb_reg = 3'b011; end
            18'b001010011011000011: begin rgb_reg = 3'b011; end
            18'b001010011011000100: begin rgb_reg = 3'b011; end
            18'b001010011011000101: begin rgb_reg = 3'b011; end
            18'b001010011011001001: begin rgb_reg = 3'b001; end
            18'b001010011011001010: begin rgb_reg = 3'b011; end
            18'b001010011011001011: begin rgb_reg = 3'b011; end
            18'b001010011011001100: begin rgb_reg = 3'b011; end
            18'b001010011011011000: begin rgb_reg = 3'b001; end
            18'b001010011011011001: begin rgb_reg = 3'b011; end
            18'b001010011011011010: begin rgb_reg = 3'b011; end
            18'b001010011011011011: begin rgb_reg = 3'b011; end
            18'b001010011011100000: begin rgb_reg = 3'b011; end
            18'b001010011011100001: begin rgb_reg = 3'b011; end
            18'b001010011011100010: begin rgb_reg = 3'b011; end
            18'b001010011011100011: begin rgb_reg = 3'b011; end
            18'b001010011011110110: begin rgb_reg = 3'b001; end
            18'b001010011011110111: begin rgb_reg = 3'b011; end
            18'b001010011011111000: begin rgb_reg = 3'b011; end
            18'b001010011011111001: begin rgb_reg = 3'b011; end
            18'b001010011100000101: begin rgb_reg = 3'b001; end
            18'b001010011100000110: begin rgb_reg = 3'b011; end
            18'b001010011100000111: begin rgb_reg = 3'b011; end
            18'b001010011100001000: begin rgb_reg = 3'b011; end
            18'b001010011100001101: begin rgb_reg = 3'b011; end
            18'b001010011100001110: begin rgb_reg = 3'b011; end
            18'b001010011100001111: begin rgb_reg = 3'b011; end
            18'b001010011100010000: begin rgb_reg = 3'b011; end
            18'b001010011100010001: begin rgb_reg = 3'b011; end
            18'b001010011100010010: begin rgb_reg = 3'b011; end
            18'b001010011100010011: begin rgb_reg = 3'b011; end
            18'b001010011100010100: begin rgb_reg = 3'b001; end
            18'b001010011100011000: begin rgb_reg = 3'b011; end
            18'b001010011100011001: begin rgb_reg = 3'b011; end
            18'b001010011100011010: begin rgb_reg = 3'b011; end
            18'b001010011100011011: begin rgb_reg = 3'b011; end
            18'b001010011100011100: begin rgb_reg = 3'b011; end
            18'b001010011100011101: begin rgb_reg = 3'b011; end
            18'b001010011100011110: begin rgb_reg = 3'b011; end
            18'b001010011100011111: begin rgb_reg = 3'b011; end
            18'b001010011100100011: begin rgb_reg = 3'b001; end
            18'b001010011100100100: begin rgb_reg = 3'b011; end
            18'b001010011100100101: begin rgb_reg = 3'b011; end
            18'b001010011100100110: begin rgb_reg = 3'b011; end
            18'b001010011100110010: begin rgb_reg = 3'b001; end
            18'b001010011100110011: begin rgb_reg = 3'b011; end
            18'b001010011100110100: begin rgb_reg = 3'b011; end
            18'b001010011100110101: begin rgb_reg = 3'b011; end
            18'b001010011100111010: begin rgb_reg = 3'b011; end
            18'b001010011100111011: begin rgb_reg = 3'b011; end
            18'b001010011100111100: begin rgb_reg = 3'b011; end
            18'b001010011100111101: begin rgb_reg = 3'b011; end
            18'b001010011101001001: begin rgb_reg = 3'b011; end
            18'b001010011101001010: begin rgb_reg = 3'b011; end
            18'b001010011101001011: begin rgb_reg = 3'b011; end
            18'b001010011101001100: begin rgb_reg = 3'b011; end
            18'b001010011101010000: begin rgb_reg = 3'b001; end
            18'b001010011101010001: begin rgb_reg = 3'b011; end
            18'b001010011101010010: begin rgb_reg = 3'b011; end
            18'b001010011101010011: begin rgb_reg = 3'b011; end
            18'b001010100010011101: begin rgb_reg = 3'b001; end
            18'b001010100010011110: begin rgb_reg = 3'b001; end
            18'b001010100010011111: begin rgb_reg = 3'b001; end
            18'b001010100010100000: begin rgb_reg = 3'b001; end
            18'b001010100010100001: begin rgb_reg = 3'b001; end
            18'b001010100010100010: begin rgb_reg = 3'b001; end
            18'b001010100010100011: begin rgb_reg = 3'b001; end
            18'b001010100010100100: begin rgb_reg = 3'b001; end
            18'b001010100010100101: begin rgb_reg = 3'b001; end
            18'b001010100010100110: begin rgb_reg = 3'b001; end
            18'b001010100010100111: begin rgb_reg = 3'b001; end
            18'b001010100010101000: begin rgb_reg = 3'b001; end
            18'b001010100010101001: begin rgb_reg = 3'b001; end
            18'b001010100010101010: begin rgb_reg = 3'b001; end
            18'b001010100010101011: begin rgb_reg = 3'b001; end
            18'b001010100010101100: begin rgb_reg = 3'b001; end
            18'b001010100010101101: begin rgb_reg = 3'b001; end
            18'b001010100010101110: begin rgb_reg = 3'b001; end
            18'b001010100010110011: begin rgb_reg = 3'b011; end
            18'b001010100010110100: begin rgb_reg = 3'b011; end
            18'b001010100010110101: begin rgb_reg = 3'b011; end
            18'b001010100010110110: begin rgb_reg = 3'b011; end
            18'b001010100011000010: begin rgb_reg = 3'b011; end
            18'b001010100011000011: begin rgb_reg = 3'b011; end
            18'b001010100011000100: begin rgb_reg = 3'b011; end
            18'b001010100011000101: begin rgb_reg = 3'b011; end
            18'b001010100011001001: begin rgb_reg = 3'b001; end
            18'b001010100011001010: begin rgb_reg = 3'b011; end
            18'b001010100011001011: begin rgb_reg = 3'b011; end
            18'b001010100011001100: begin rgb_reg = 3'b011; end
            18'b001010100011001101: begin rgb_reg = 3'b001; end
            18'b001010100011001110: begin rgb_reg = 3'b001; end
            18'b001010100011001111: begin rgb_reg = 3'b001; end
            18'b001010100011010000: begin rgb_reg = 3'b001; end
            18'b001010100011010001: begin rgb_reg = 3'b001; end
            18'b001010100011010010: begin rgb_reg = 3'b001; end
            18'b001010100011010011: begin rgb_reg = 3'b001; end
            18'b001010100011010100: begin rgb_reg = 3'b001; end
            18'b001010100011010101: begin rgb_reg = 3'b001; end
            18'b001010100011010110: begin rgb_reg = 3'b001; end
            18'b001010100011010111: begin rgb_reg = 3'b001; end
            18'b001010100011011000: begin rgb_reg = 3'b001; end
            18'b001010100011011001: begin rgb_reg = 3'b001; end
            18'b001010100011011010: begin rgb_reg = 3'b001; end
            18'b001010100011011011: begin rgb_reg = 3'b001; end
            18'b001010100011100000: begin rgb_reg = 3'b011; end
            18'b001010100011100001: begin rgb_reg = 3'b011; end
            18'b001010100011100010: begin rgb_reg = 3'b011; end
            18'b001010100011100011: begin rgb_reg = 3'b011; end
            18'b001010100011100100: begin rgb_reg = 3'b001; end
            18'b001010100011100101: begin rgb_reg = 3'b001; end
            18'b001010100011100110: begin rgb_reg = 3'b001; end
            18'b001010100011100111: begin rgb_reg = 3'b001; end
            18'b001010100011101000: begin rgb_reg = 3'b001; end
            18'b001010100011101001: begin rgb_reg = 3'b001; end
            18'b001010100011101010: begin rgb_reg = 3'b001; end
            18'b001010100011101011: begin rgb_reg = 3'b001; end
            18'b001010100011101100: begin rgb_reg = 3'b001; end
            18'b001010100011101101: begin rgb_reg = 3'b001; end
            18'b001010100011101110: begin rgb_reg = 3'b001; end
            18'b001010100011101111: begin rgb_reg = 3'b001; end
            18'b001010100011110000: begin rgb_reg = 3'b001; end
            18'b001010100011110001: begin rgb_reg = 3'b001; end
            18'b001010100011110010: begin rgb_reg = 3'b001; end
            18'b001010100011110110: begin rgb_reg = 3'b001; end
            18'b001010100011110111: begin rgb_reg = 3'b011; end
            18'b001010100011111000: begin rgb_reg = 3'b011; end
            18'b001010100011111001: begin rgb_reg = 3'b011; end
            18'b001010100100000101: begin rgb_reg = 3'b001; end
            18'b001010100100000110: begin rgb_reg = 3'b011; end
            18'b001010100100000111: begin rgb_reg = 3'b011; end
            18'b001010100100001000: begin rgb_reg = 3'b011; end
            18'b001010100100001101: begin rgb_reg = 3'b011; end
            18'b001010100100001110: begin rgb_reg = 3'b011; end
            18'b001010100100001111: begin rgb_reg = 3'b011; end
            18'b001010100100010000: begin rgb_reg = 3'b011; end
            18'b001010100100010001: begin rgb_reg = 3'b001; end
            18'b001010100100010010: begin rgb_reg = 3'b001; end
            18'b001010100100010011: begin rgb_reg = 3'b001; end
            18'b001010100100011000: begin rgb_reg = 3'b001; end
            18'b001010100100011001: begin rgb_reg = 3'b001; end
            18'b001010100100011010: begin rgb_reg = 3'b001; end
            18'b001010100100011011: begin rgb_reg = 3'b001; end
            18'b001010100100011100: begin rgb_reg = 3'b011; end
            18'b001010100100011101: begin rgb_reg = 3'b011; end
            18'b001010100100011110: begin rgb_reg = 3'b011; end
            18'b001010100100011111: begin rgb_reg = 3'b011; end
            18'b001010100100100011: begin rgb_reg = 3'b001; end
            18'b001010100100100100: begin rgb_reg = 3'b011; end
            18'b001010100100100101: begin rgb_reg = 3'b011; end
            18'b001010100100100110: begin rgb_reg = 3'b011; end
            18'b001010100100110010: begin rgb_reg = 3'b001; end
            18'b001010100100110011: begin rgb_reg = 3'b011; end
            18'b001010100100110100: begin rgb_reg = 3'b011; end
            18'b001010100100110101: begin rgb_reg = 3'b011; end
            18'b001010100100111010: begin rgb_reg = 3'b011; end
            18'b001010100100111011: begin rgb_reg = 3'b011; end
            18'b001010100100111100: begin rgb_reg = 3'b011; end
            18'b001010100100111101: begin rgb_reg = 3'b011; end
            18'b001010100101001001: begin rgb_reg = 3'b011; end
            18'b001010100101001010: begin rgb_reg = 3'b011; end
            18'b001010100101001011: begin rgb_reg = 3'b011; end
            18'b001010100101001100: begin rgb_reg = 3'b011; end
            18'b001010100101010000: begin rgb_reg = 3'b001; end
            18'b001010100101010001: begin rgb_reg = 3'b011; end
            18'b001010100101010010: begin rgb_reg = 3'b011; end
            18'b001010100101010011: begin rgb_reg = 3'b011; end
            18'b001010100101010100: begin rgb_reg = 3'b001; end
            18'b001010100101010101: begin rgb_reg = 3'b001; end
            18'b001010100101010110: begin rgb_reg = 3'b001; end
            18'b001010100101010111: begin rgb_reg = 3'b001; end
            18'b001010100101011000: begin rgb_reg = 3'b001; end
            18'b001010100101011001: begin rgb_reg = 3'b001; end
            18'b001010100101011010: begin rgb_reg = 3'b001; end
            18'b001010100101011011: begin rgb_reg = 3'b001; end
            18'b001010100101011100: begin rgb_reg = 3'b001; end
            18'b001010100101011101: begin rgb_reg = 3'b001; end
            18'b001010100101011110: begin rgb_reg = 3'b001; end
            18'b001010100101011111: begin rgb_reg = 3'b001; end
            18'b001010100101100000: begin rgb_reg = 3'b001; end
            18'b001010100101100001: begin rgb_reg = 3'b001; end
            18'b001010100101100010: begin rgb_reg = 3'b001; end
            18'b001010101010100000: begin rgb_reg = 3'b011; end
            18'b001010101010100001: begin rgb_reg = 3'b011; end
            18'b001010101010100010: begin rgb_reg = 3'b011; end
            18'b001010101010100011: begin rgb_reg = 3'b011; end
            18'b001010101010100100: begin rgb_reg = 3'b011; end
            18'b001010101010100101: begin rgb_reg = 3'b011; end
            18'b001010101010100110: begin rgb_reg = 3'b011; end
            18'b001010101010100111: begin rgb_reg = 3'b011; end
            18'b001010101010101000: begin rgb_reg = 3'b011; end
            18'b001010101010101001: begin rgb_reg = 3'b011; end
            18'b001010101010101010: begin rgb_reg = 3'b011; end
            18'b001010101010101011: begin rgb_reg = 3'b001; end
            18'b001010101010110011: begin rgb_reg = 3'b011; end
            18'b001010101010110100: begin rgb_reg = 3'b011; end
            18'b001010101010110101: begin rgb_reg = 3'b011; end
            18'b001010101010110110: begin rgb_reg = 3'b011; end
            18'b001010101011000010: begin rgb_reg = 3'b011; end
            18'b001010101011000011: begin rgb_reg = 3'b011; end
            18'b001010101011000100: begin rgb_reg = 3'b011; end
            18'b001010101011000101: begin rgb_reg = 3'b011; end
            18'b001010101011001001: begin rgb_reg = 3'b001; end
            18'b001010101011001010: begin rgb_reg = 3'b011; end
            18'b001010101011001011: begin rgb_reg = 3'b011; end
            18'b001010101011001100: begin rgb_reg = 3'b011; end
            18'b001010101011001101: begin rgb_reg = 3'b011; end
            18'b001010101011001110: begin rgb_reg = 3'b011; end
            18'b001010101011001111: begin rgb_reg = 3'b011; end
            18'b001010101011010000: begin rgb_reg = 3'b011; end
            18'b001010101011010001: begin rgb_reg = 3'b011; end
            18'b001010101011010010: begin rgb_reg = 3'b011; end
            18'b001010101011010011: begin rgb_reg = 3'b011; end
            18'b001010101011010100: begin rgb_reg = 3'b011; end
            18'b001010101011010101: begin rgb_reg = 3'b011; end
            18'b001010101011010110: begin rgb_reg = 3'b011; end
            18'b001010101011010111: begin rgb_reg = 3'b011; end
            18'b001010101011011000: begin rgb_reg = 3'b001; end
            18'b001010101011100000: begin rgb_reg = 3'b011; end
            18'b001010101011100001: begin rgb_reg = 3'b011; end
            18'b001010101011100010: begin rgb_reg = 3'b011; end
            18'b001010101011100011: begin rgb_reg = 3'b011; end
            18'b001010101011100100: begin rgb_reg = 3'b011; end
            18'b001010101011100101: begin rgb_reg = 3'b011; end
            18'b001010101011100110: begin rgb_reg = 3'b011; end
            18'b001010101011100111: begin rgb_reg = 3'b011; end
            18'b001010101011101000: begin rgb_reg = 3'b011; end
            18'b001010101011101001: begin rgb_reg = 3'b011; end
            18'b001010101011101010: begin rgb_reg = 3'b011; end
            18'b001010101011101011: begin rgb_reg = 3'b011; end
            18'b001010101011101100: begin rgb_reg = 3'b011; end
            18'b001010101011101101: begin rgb_reg = 3'b011; end
            18'b001010101011101110: begin rgb_reg = 3'b011; end
            18'b001010101011101111: begin rgb_reg = 3'b011; end
            18'b001010101011110000: begin rgb_reg = 3'b011; end
            18'b001010101011110001: begin rgb_reg = 3'b011; end
            18'b001010101011110010: begin rgb_reg = 3'b011; end
            18'b001010101011110110: begin rgb_reg = 3'b001; end
            18'b001010101011110111: begin rgb_reg = 3'b011; end
            18'b001010101011111000: begin rgb_reg = 3'b011; end
            18'b001010101011111001: begin rgb_reg = 3'b011; end
            18'b001010101100000101: begin rgb_reg = 3'b001; end
            18'b001010101100000110: begin rgb_reg = 3'b011; end
            18'b001010101100000111: begin rgb_reg = 3'b011; end
            18'b001010101100001000: begin rgb_reg = 3'b011; end
            18'b001010101100001101: begin rgb_reg = 3'b011; end
            18'b001010101100001110: begin rgb_reg = 3'b011; end
            18'b001010101100001111: begin rgb_reg = 3'b011; end
            18'b001010101100010000: begin rgb_reg = 3'b011; end
            18'b001010101100011100: begin rgb_reg = 3'b011; end
            18'b001010101100011101: begin rgb_reg = 3'b011; end
            18'b001010101100011110: begin rgb_reg = 3'b011; end
            18'b001010101100011111: begin rgb_reg = 3'b011; end
            18'b001010101100100011: begin rgb_reg = 3'b001; end
            18'b001010101100100100: begin rgb_reg = 3'b011; end
            18'b001010101100100101: begin rgb_reg = 3'b011; end
            18'b001010101100100110: begin rgb_reg = 3'b011; end
            18'b001010101100110010: begin rgb_reg = 3'b001; end
            18'b001010101100110011: begin rgb_reg = 3'b011; end
            18'b001010101100110100: begin rgb_reg = 3'b011; end
            18'b001010101100110101: begin rgb_reg = 3'b011; end
            18'b001010101100111010: begin rgb_reg = 3'b011; end
            18'b001010101100111011: begin rgb_reg = 3'b011; end
            18'b001010101100111100: begin rgb_reg = 3'b011; end
            18'b001010101100111101: begin rgb_reg = 3'b011; end
            18'b001010101101001001: begin rgb_reg = 3'b011; end
            18'b001010101101001010: begin rgb_reg = 3'b011; end
            18'b001010101101001011: begin rgb_reg = 3'b011; end
            18'b001010101101001100: begin rgb_reg = 3'b011; end
            18'b001010101101010000: begin rgb_reg = 3'b001; end
            18'b001010101101010001: begin rgb_reg = 3'b011; end
            18'b001010101101010010: begin rgb_reg = 3'b011; end
            18'b001010101101010011: begin rgb_reg = 3'b011; end
            18'b001010101101010100: begin rgb_reg = 3'b011; end
            18'b001010101101010101: begin rgb_reg = 3'b011; end
            18'b001010101101010110: begin rgb_reg = 3'b011; end
            18'b001010101101010111: begin rgb_reg = 3'b011; end
            18'b001010101101011000: begin rgb_reg = 3'b011; end
            18'b001010101101011001: begin rgb_reg = 3'b011; end
            18'b001010101101011010: begin rgb_reg = 3'b011; end
            18'b001010101101011011: begin rgb_reg = 3'b011; end
            18'b001010101101011100: begin rgb_reg = 3'b011; end
            18'b001010101101011101: begin rgb_reg = 3'b011; end
            18'b001010101101011110: begin rgb_reg = 3'b011; end
            18'b001010101101011111: begin rgb_reg = 3'b011; end
            18'b001010101101100000: begin rgb_reg = 3'b011; end
            18'b001010101101100001: begin rgb_reg = 3'b011; end
            18'b001010101101100010: begin rgb_reg = 3'b011; end
            18'b001010110010100000: begin rgb_reg = 3'b011; end
            18'b001010110010100001: begin rgb_reg = 3'b011; end
            18'b001010110010100010: begin rgb_reg = 3'b011; end
            18'b001010110010100011: begin rgb_reg = 3'b011; end
            18'b001010110010100100: begin rgb_reg = 3'b011; end
            18'b001010110010100101: begin rgb_reg = 3'b011; end
            18'b001010110010100110: begin rgb_reg = 3'b011; end
            18'b001010110010100111: begin rgb_reg = 3'b011; end
            18'b001010110010101000: begin rgb_reg = 3'b011; end
            18'b001010110010101001: begin rgb_reg = 3'b011; end
            18'b001010110010101010: begin rgb_reg = 3'b011; end
            18'b001010110010101011: begin rgb_reg = 3'b001; end
            18'b001010110010110011: begin rgb_reg = 3'b011; end
            18'b001010110010110100: begin rgb_reg = 3'b011; end
            18'b001010110010110101: begin rgb_reg = 3'b011; end
            18'b001010110010110110: begin rgb_reg = 3'b011; end
            18'b001010110011000010: begin rgb_reg = 3'b011; end
            18'b001010110011000011: begin rgb_reg = 3'b011; end
            18'b001010110011000100: begin rgb_reg = 3'b011; end
            18'b001010110011000101: begin rgb_reg = 3'b011; end
            18'b001010110011001001: begin rgb_reg = 3'b001; end
            18'b001010110011001010: begin rgb_reg = 3'b011; end
            18'b001010110011001011: begin rgb_reg = 3'b011; end
            18'b001010110011001100: begin rgb_reg = 3'b011; end
            18'b001010110011001101: begin rgb_reg = 3'b011; end
            18'b001010110011001110: begin rgb_reg = 3'b011; end
            18'b001010110011001111: begin rgb_reg = 3'b011; end
            18'b001010110011010000: begin rgb_reg = 3'b011; end
            18'b001010110011010001: begin rgb_reg = 3'b011; end
            18'b001010110011010010: begin rgb_reg = 3'b011; end
            18'b001010110011010011: begin rgb_reg = 3'b011; end
            18'b001010110011010100: begin rgb_reg = 3'b011; end
            18'b001010110011010101: begin rgb_reg = 3'b011; end
            18'b001010110011010110: begin rgb_reg = 3'b011; end
            18'b001010110011010111: begin rgb_reg = 3'b011; end
            18'b001010110011011000: begin rgb_reg = 3'b001; end
            18'b001010110011100000: begin rgb_reg = 3'b011; end
            18'b001010110011100001: begin rgb_reg = 3'b011; end
            18'b001010110011100010: begin rgb_reg = 3'b011; end
            18'b001010110011100011: begin rgb_reg = 3'b011; end
            18'b001010110011100100: begin rgb_reg = 3'b011; end
            18'b001010110011100101: begin rgb_reg = 3'b011; end
            18'b001010110011100110: begin rgb_reg = 3'b011; end
            18'b001010110011100111: begin rgb_reg = 3'b011; end
            18'b001010110011101000: begin rgb_reg = 3'b011; end
            18'b001010110011101001: begin rgb_reg = 3'b011; end
            18'b001010110011101010: begin rgb_reg = 3'b011; end
            18'b001010110011101011: begin rgb_reg = 3'b011; end
            18'b001010110011101100: begin rgb_reg = 3'b011; end
            18'b001010110011101101: begin rgb_reg = 3'b011; end
            18'b001010110011101110: begin rgb_reg = 3'b011; end
            18'b001010110011101111: begin rgb_reg = 3'b011; end
            18'b001010110011110000: begin rgb_reg = 3'b011; end
            18'b001010110011110001: begin rgb_reg = 3'b011; end
            18'b001010110011110010: begin rgb_reg = 3'b011; end
            18'b001010110011110110: begin rgb_reg = 3'b001; end
            18'b001010110011110111: begin rgb_reg = 3'b011; end
            18'b001010110011111000: begin rgb_reg = 3'b011; end
            18'b001010110011111001: begin rgb_reg = 3'b011; end
            18'b001010110100000101: begin rgb_reg = 3'b001; end
            18'b001010110100000110: begin rgb_reg = 3'b011; end
            18'b001010110100000111: begin rgb_reg = 3'b011; end
            18'b001010110100001000: begin rgb_reg = 3'b011; end
            18'b001010110100001101: begin rgb_reg = 3'b011; end
            18'b001010110100001110: begin rgb_reg = 3'b011; end
            18'b001010110100001111: begin rgb_reg = 3'b011; end
            18'b001010110100010000: begin rgb_reg = 3'b011; end
            18'b001010110100011100: begin rgb_reg = 3'b011; end
            18'b001010110100011101: begin rgb_reg = 3'b011; end
            18'b001010110100011110: begin rgb_reg = 3'b011; end
            18'b001010110100011111: begin rgb_reg = 3'b011; end
            18'b001010110100100011: begin rgb_reg = 3'b001; end
            18'b001010110100100100: begin rgb_reg = 3'b011; end
            18'b001010110100100101: begin rgb_reg = 3'b011; end
            18'b001010110100100110: begin rgb_reg = 3'b011; end
            18'b001010110100110010: begin rgb_reg = 3'b001; end
            18'b001010110100110011: begin rgb_reg = 3'b011; end
            18'b001010110100110100: begin rgb_reg = 3'b011; end
            18'b001010110100110101: begin rgb_reg = 3'b011; end
            18'b001010110100111010: begin rgb_reg = 3'b011; end
            18'b001010110100111011: begin rgb_reg = 3'b011; end
            18'b001010110100111100: begin rgb_reg = 3'b011; end
            18'b001010110100111101: begin rgb_reg = 3'b011; end
            18'b001010110101001001: begin rgb_reg = 3'b011; end
            18'b001010110101001010: begin rgb_reg = 3'b011; end
            18'b001010110101001011: begin rgb_reg = 3'b011; end
            18'b001010110101001100: begin rgb_reg = 3'b011; end
            18'b001010110101010000: begin rgb_reg = 3'b001; end
            18'b001010110101010001: begin rgb_reg = 3'b011; end
            18'b001010110101010010: begin rgb_reg = 3'b011; end
            18'b001010110101010011: begin rgb_reg = 3'b011; end
            18'b001010110101010100: begin rgb_reg = 3'b011; end
            18'b001010110101010101: begin rgb_reg = 3'b011; end
            18'b001010110101010110: begin rgb_reg = 3'b011; end
            18'b001010110101010111: begin rgb_reg = 3'b011; end
            18'b001010110101011000: begin rgb_reg = 3'b011; end
            18'b001010110101011001: begin rgb_reg = 3'b011; end
            18'b001010110101011010: begin rgb_reg = 3'b011; end
            18'b001010110101011011: begin rgb_reg = 3'b011; end
            18'b001010110101011100: begin rgb_reg = 3'b011; end
            18'b001010110101011101: begin rgb_reg = 3'b011; end
            18'b001010110101011110: begin rgb_reg = 3'b011; end
            18'b001010110101011111: begin rgb_reg = 3'b011; end
            18'b001010110101100000: begin rgb_reg = 3'b011; end
            18'b001010110101100001: begin rgb_reg = 3'b011; end
            18'b001010110101100010: begin rgb_reg = 3'b011; end
            18'b001010111010100000: begin rgb_reg = 3'b011; end
            18'b001010111010100001: begin rgb_reg = 3'b011; end
            18'b001010111010100010: begin rgb_reg = 3'b011; end
            18'b001010111010100011: begin rgb_reg = 3'b011; end
            18'b001010111010100100: begin rgb_reg = 3'b011; end
            18'b001010111010100101: begin rgb_reg = 3'b011; end
            18'b001010111010100110: begin rgb_reg = 3'b011; end
            18'b001010111010100111: begin rgb_reg = 3'b011; end
            18'b001010111010101000: begin rgb_reg = 3'b011; end
            18'b001010111010101001: begin rgb_reg = 3'b011; end
            18'b001010111010101010: begin rgb_reg = 3'b011; end
            18'b001010111010101011: begin rgb_reg = 3'b001; end
            18'b001010111010110011: begin rgb_reg = 3'b011; end
            18'b001010111010110100: begin rgb_reg = 3'b011; end
            18'b001010111010110101: begin rgb_reg = 3'b011; end
            18'b001010111010110110: begin rgb_reg = 3'b011; end
            18'b001010111011000010: begin rgb_reg = 3'b011; end
            18'b001010111011000011: begin rgb_reg = 3'b011; end
            18'b001010111011000100: begin rgb_reg = 3'b011; end
            18'b001010111011000101: begin rgb_reg = 3'b011; end
            18'b001010111011001001: begin rgb_reg = 3'b001; end
            18'b001010111011001010: begin rgb_reg = 3'b011; end
            18'b001010111011001011: begin rgb_reg = 3'b011; end
            18'b001010111011001100: begin rgb_reg = 3'b011; end
            18'b001010111011001101: begin rgb_reg = 3'b011; end
            18'b001010111011001110: begin rgb_reg = 3'b011; end
            18'b001010111011001111: begin rgb_reg = 3'b011; end
            18'b001010111011010000: begin rgb_reg = 3'b011; end
            18'b001010111011010001: begin rgb_reg = 3'b011; end
            18'b001010111011010010: begin rgb_reg = 3'b011; end
            18'b001010111011010011: begin rgb_reg = 3'b011; end
            18'b001010111011010100: begin rgb_reg = 3'b011; end
            18'b001010111011010101: begin rgb_reg = 3'b011; end
            18'b001010111011010110: begin rgb_reg = 3'b011; end
            18'b001010111011010111: begin rgb_reg = 3'b011; end
            18'b001010111011011000: begin rgb_reg = 3'b001; end
            18'b001010111011100000: begin rgb_reg = 3'b011; end
            18'b001010111011100001: begin rgb_reg = 3'b011; end
            18'b001010111011100010: begin rgb_reg = 3'b011; end
            18'b001010111011100011: begin rgb_reg = 3'b011; end
            18'b001010111011100100: begin rgb_reg = 3'b011; end
            18'b001010111011100101: begin rgb_reg = 3'b011; end
            18'b001010111011100110: begin rgb_reg = 3'b011; end
            18'b001010111011100111: begin rgb_reg = 3'b011; end
            18'b001010111011101000: begin rgb_reg = 3'b011; end
            18'b001010111011101001: begin rgb_reg = 3'b011; end
            18'b001010111011101010: begin rgb_reg = 3'b011; end
            18'b001010111011101011: begin rgb_reg = 3'b011; end
            18'b001010111011101100: begin rgb_reg = 3'b011; end
            18'b001010111011101101: begin rgb_reg = 3'b011; end
            18'b001010111011101110: begin rgb_reg = 3'b011; end
            18'b001010111011101111: begin rgb_reg = 3'b011; end
            18'b001010111011110000: begin rgb_reg = 3'b011; end
            18'b001010111011110001: begin rgb_reg = 3'b011; end
            18'b001010111011110010: begin rgb_reg = 3'b011; end
            18'b001010111011110110: begin rgb_reg = 3'b001; end
            18'b001010111011110111: begin rgb_reg = 3'b011; end
            18'b001010111011111000: begin rgb_reg = 3'b011; end
            18'b001010111011111001: begin rgb_reg = 3'b011; end
            18'b001010111100000101: begin rgb_reg = 3'b001; end
            18'b001010111100000110: begin rgb_reg = 3'b011; end
            18'b001010111100000111: begin rgb_reg = 3'b011; end
            18'b001010111100001000: begin rgb_reg = 3'b011; end
            18'b001010111100001101: begin rgb_reg = 3'b011; end
            18'b001010111100001110: begin rgb_reg = 3'b011; end
            18'b001010111100001111: begin rgb_reg = 3'b011; end
            18'b001010111100010000: begin rgb_reg = 3'b011; end
            18'b001010111100011100: begin rgb_reg = 3'b011; end
            18'b001010111100011101: begin rgb_reg = 3'b011; end
            18'b001010111100011110: begin rgb_reg = 3'b011; end
            18'b001010111100011111: begin rgb_reg = 3'b011; end
            18'b001010111100100011: begin rgb_reg = 3'b001; end
            18'b001010111100100100: begin rgb_reg = 3'b011; end
            18'b001010111100100101: begin rgb_reg = 3'b011; end
            18'b001010111100100110: begin rgb_reg = 3'b011; end
            18'b001010111100110010: begin rgb_reg = 3'b001; end
            18'b001010111100110011: begin rgb_reg = 3'b011; end
            18'b001010111100110100: begin rgb_reg = 3'b011; end
            18'b001010111100110101: begin rgb_reg = 3'b011; end
            18'b001010111100111010: begin rgb_reg = 3'b011; end
            18'b001010111100111011: begin rgb_reg = 3'b011; end
            18'b001010111100111100: begin rgb_reg = 3'b011; end
            18'b001010111100111101: begin rgb_reg = 3'b011; end
            18'b001010111101001001: begin rgb_reg = 3'b011; end
            18'b001010111101001010: begin rgb_reg = 3'b011; end
            18'b001010111101001011: begin rgb_reg = 3'b011; end
            18'b001010111101001100: begin rgb_reg = 3'b011; end
            18'b001010111101010000: begin rgb_reg = 3'b001; end
            18'b001010111101010001: begin rgb_reg = 3'b011; end
            18'b001010111101010010: begin rgb_reg = 3'b011; end
            18'b001010111101010011: begin rgb_reg = 3'b011; end
            18'b001010111101010100: begin rgb_reg = 3'b011; end
            18'b001010111101010101: begin rgb_reg = 3'b011; end
            18'b001010111101010110: begin rgb_reg = 3'b011; end
            18'b001010111101010111: begin rgb_reg = 3'b011; end
            18'b001010111101011000: begin rgb_reg = 3'b011; end
            18'b001010111101011001: begin rgb_reg = 3'b011; end
            18'b001010111101011010: begin rgb_reg = 3'b011; end
            18'b001010111101011011: begin rgb_reg = 3'b011; end
            18'b001010111101011100: begin rgb_reg = 3'b011; end
            18'b001010111101011101: begin rgb_reg = 3'b011; end
            18'b001010111101011110: begin rgb_reg = 3'b011; end
            18'b001010111101011111: begin rgb_reg = 3'b011; end
            18'b001010111101100000: begin rgb_reg = 3'b011; end
            18'b001010111101100001: begin rgb_reg = 3'b011; end
            18'b001010111101100010: begin rgb_reg = 3'b011; end
            18'b001110011011110110: begin rgb_reg = 3'b111; end
            18'b001110011011110111: begin rgb_reg = 3'b111; end
            18'b001110100011110110: begin rgb_reg = 3'b111; end
            18'b001110100011110111: begin rgb_reg = 3'b111; end
            18'b001110101011110110: begin rgb_reg = 3'b111; end
            18'b001110101011110111: begin rgb_reg = 3'b111; end
            18'b001110110011110110: begin rgb_reg = 3'b111; end
            18'b001110110011110111: begin rgb_reg = 3'b111; end
            18'b001110111011110110: begin rgb_reg = 3'b111; end
            18'b001110111011110111: begin rgb_reg = 3'b111; end
            18'b001110111011111010: begin rgb_reg = 3'b111; end
            18'b001110111011111011: begin rgb_reg = 3'b111; end
            18'b001110111011111100: begin rgb_reg = 3'b111; end
            18'b001110111100000001: begin rgb_reg = 3'b111; end
            18'b001110111100001000: begin rgb_reg = 3'b111; end
            18'b001111000011110110: begin rgb_reg = 3'b111; end
            18'b001111000011110111: begin rgb_reg = 3'b111; end
            18'b001111000011111000: begin rgb_reg = 3'b111; end
            18'b001111000011111101: begin rgb_reg = 3'b111; end
            18'b001111000100000001: begin rgb_reg = 3'b111; end
            18'b001111000100001000: begin rgb_reg = 3'b111; end
            18'b001111001011110110: begin rgb_reg = 3'b111; end
            18'b001111001011110111: begin rgb_reg = 3'b111; end
            18'b001111001011111000: begin rgb_reg = 3'b111; end
            18'b001111001011111101: begin rgb_reg = 3'b111; end
            18'b001111001011111110: begin rgb_reg = 3'b111; end
            18'b001111001100000001: begin rgb_reg = 3'b111; end
            18'b001111001100001000: begin rgb_reg = 3'b111; end
            18'b001111010011110110: begin rgb_reg = 3'b111; end
            18'b001111010011110111: begin rgb_reg = 3'b111; end
            18'b001111010011111101: begin rgb_reg = 3'b111; end
            18'b001111010011111110: begin rgb_reg = 3'b111; end
            18'b001111010100000001: begin rgb_reg = 3'b111; end
            18'b001111010100001000: begin rgb_reg = 3'b111; end
            18'b001111011011110110: begin rgb_reg = 3'b111; end
            18'b001111011011110111: begin rgb_reg = 3'b111; end
            18'b001111011011111101: begin rgb_reg = 3'b111; end
            18'b001111011011111110: begin rgb_reg = 3'b111; end
            18'b001111011100000001: begin rgb_reg = 3'b111; end
            18'b001111011100001000: begin rgb_reg = 3'b111; end
            18'b001111100011110110: begin rgb_reg = 3'b111; end
            18'b001111100011110111: begin rgb_reg = 3'b111; end
            18'b001111100011111101: begin rgb_reg = 3'b111; end
            18'b001111100011111110: begin rgb_reg = 3'b111; end
            18'b001111100100000010: begin rgb_reg = 3'b111; end
            18'b001111100100000011: begin rgb_reg = 3'b111; end
            18'b001111100100000100: begin rgb_reg = 3'b111; end
            18'b001111100100000101: begin rgb_reg = 3'b111; end
            18'b001111100100000110: begin rgb_reg = 3'b111; end
            18'b001111100100000111: begin rgb_reg = 3'b111; end
            18'b001111100100001000: begin rgb_reg = 3'b111; end
            18'b001111101011110110: begin rgb_reg = 3'b111; end
            18'b001111101011110111: begin rgb_reg = 3'b111; end
            18'b001111101100000111: begin rgb_reg = 3'b111; end
            18'b001111101100001000: begin rgb_reg = 3'b111; end
            18'b001111110011110110: begin rgb_reg = 3'b111; end
            18'b001111110011110111: begin rgb_reg = 3'b111; end
            18'b001111110011111000: begin rgb_reg = 3'b111; end
            18'b001111110011111001: begin rgb_reg = 3'b111; end
            18'b001111110011111010: begin rgb_reg = 3'b111; end
            18'b001111110011111011: begin rgb_reg = 3'b111; end
            18'b001111110011111100: begin rgb_reg = 3'b111; end
            18'b001111110100001000: begin rgb_reg = 3'b111; end
            18'b001111111100000001: begin rgb_reg = 3'b111; end
            18'b001111111100000010: begin rgb_reg = 3'b111; end
            18'b001111111100000011: begin rgb_reg = 3'b111; end
            18'b001111111100000100: begin rgb_reg = 3'b111; end
            18'b001111111100000101: begin rgb_reg = 3'b111; end
            18'b001111111100000110: begin rgb_reg = 3'b111; end
            18'b010000000100000001: begin rgb_reg = 3'b111; end
            18'b010000000100000010: begin rgb_reg = 3'b111; end
            18'b010000000100000011: begin rgb_reg = 3'b111; end
            18'b010000000100000100: begin rgb_reg = 3'b111; end
            18'b010000000100000101: begin rgb_reg = 3'b111; end
            18'b010000000100000110: begin rgb_reg = 3'b111; end
            18'b010010010011000010: begin rgb_reg = 3'b111; end
            18'b010010010011000011: begin rgb_reg = 3'b111; end
            18'b010010010011000100: begin rgb_reg = 3'b111; end
            18'b010010010011000101: begin rgb_reg = 3'b111; end
            18'b010010010011000110: begin rgb_reg = 3'b111; end
            18'b010010010011001101: begin rgb_reg = 3'b111; end
            18'b010010010011001110: begin rgb_reg = 3'b111; end
            18'b010010010011001111: begin rgb_reg = 3'b111; end
            18'b010010010011010000: begin rgb_reg = 3'b111; end
            18'b010010010011010001: begin rgb_reg = 3'b111; end
            18'b010010010011010010: begin rgb_reg = 3'b111; end
            18'b010010010011010011: begin rgb_reg = 3'b111; end
            18'b010010010011011011: begin rgb_reg = 3'b111; end
            18'b010010010011011100: begin rgb_reg = 3'b111; end
            18'b010010010011011101: begin rgb_reg = 3'b111; end
            18'b010010010011011110: begin rgb_reg = 3'b111; end
            18'b010010010011011111: begin rgb_reg = 3'b111; end
            18'b010010010011100000: begin rgb_reg = 3'b111; end
            18'b010010010011100001: begin rgb_reg = 3'b111; end
            18'b010010010011101011: begin rgb_reg = 3'b111; end
            18'b010010010011101100: begin rgb_reg = 3'b111; end
            18'b010010010011110110: begin rgb_reg = 3'b111; end
            18'b010010010011110111: begin rgb_reg = 3'b111; end
            18'b010010010011111000: begin rgb_reg = 3'b111; end
            18'b010010010011111001: begin rgb_reg = 3'b111; end
            18'b010010010011111010: begin rgb_reg = 3'b111; end
            18'b010010010011111011: begin rgb_reg = 3'b111; end
            18'b010010010011111100: begin rgb_reg = 3'b111; end
            18'b010010010100000001: begin rgb_reg = 3'b111; end
            18'b010010010100000010: begin rgb_reg = 3'b111; end
            18'b010010010100000011: begin rgb_reg = 3'b111; end
            18'b010010010100000100: begin rgb_reg = 3'b111; end
            18'b010010010100000101: begin rgb_reg = 3'b111; end
            18'b010010010100000110: begin rgb_reg = 3'b111; end
            18'b010010010100000111: begin rgb_reg = 3'b111; end
            18'b010010010100001000: begin rgb_reg = 3'b111; end
            18'b010010010100001001: begin rgb_reg = 3'b111; end
            18'b010010010100001010: begin rgb_reg = 3'b111; end
            18'b010010010100001011: begin rgb_reg = 3'b111; end
            18'b010010010100001100: begin rgb_reg = 3'b111; end
            18'b010010010100010011: begin rgb_reg = 3'b111; end
            18'b010010010100010100: begin rgb_reg = 3'b111; end
            18'b010010010100010101: begin rgb_reg = 3'b111; end
            18'b010010010100011110: begin rgb_reg = 3'b111; end
            18'b010010010100011111: begin rgb_reg = 3'b111; end
            18'b010010010100100000: begin rgb_reg = 3'b111; end
            18'b010010010100100001: begin rgb_reg = 3'b111; end
            18'b010010010100100010: begin rgb_reg = 3'b111; end
            18'b010010010100100011: begin rgb_reg = 3'b111; end
            18'b010010010100100100: begin rgb_reg = 3'b111; end
            18'b010010010100101100: begin rgb_reg = 3'b111; end
            18'b010010010100101101: begin rgb_reg = 3'b111; end
            18'b010010010100101110: begin rgb_reg = 3'b111; end
            18'b010010010100101111: begin rgb_reg = 3'b111; end
            18'b010010010100110000: begin rgb_reg = 3'b111; end
            18'b010010010100110001: begin rgb_reg = 3'b111; end
            18'b010010010100110010: begin rgb_reg = 3'b111; end
            18'b010010010100111100: begin rgb_reg = 3'b111; end
            18'b010010010100111101: begin rgb_reg = 3'b111; end
            18'b010010011011000010: begin rgb_reg = 3'b111; end
            18'b010010011011000011: begin rgb_reg = 3'b111; end
            18'b010010011011000100: begin rgb_reg = 3'b111; end
            18'b010010011011000101: begin rgb_reg = 3'b111; end
            18'b010010011011000110: begin rgb_reg = 3'b111; end
            18'b010010011011001101: begin rgb_reg = 3'b111; end
            18'b010010011011001110: begin rgb_reg = 3'b111; end
            18'b010010011011001111: begin rgb_reg = 3'b111; end
            18'b010010011011010000: begin rgb_reg = 3'b111; end
            18'b010010011011010001: begin rgb_reg = 3'b111; end
            18'b010010011011010010: begin rgb_reg = 3'b111; end
            18'b010010011011010011: begin rgb_reg = 3'b111; end
            18'b010010011011011011: begin rgb_reg = 3'b111; end
            18'b010010011011011100: begin rgb_reg = 3'b111; end
            18'b010010011011011101: begin rgb_reg = 3'b111; end
            18'b010010011011011110: begin rgb_reg = 3'b111; end
            18'b010010011011011111: begin rgb_reg = 3'b111; end
            18'b010010011011100000: begin rgb_reg = 3'b111; end
            18'b010010011011100001: begin rgb_reg = 3'b111; end
            18'b010010011011101011: begin rgb_reg = 3'b111; end
            18'b010010011011101100: begin rgb_reg = 3'b111; end
            18'b010010011011110110: begin rgb_reg = 3'b111; end
            18'b010010011011110111: begin rgb_reg = 3'b111; end
            18'b010010011011111000: begin rgb_reg = 3'b111; end
            18'b010010011011111001: begin rgb_reg = 3'b111; end
            18'b010010011011111010: begin rgb_reg = 3'b111; end
            18'b010010011011111011: begin rgb_reg = 3'b111; end
            18'b010010011011111100: begin rgb_reg = 3'b111; end
            18'b010010011100000001: begin rgb_reg = 3'b111; end
            18'b010010011100000010: begin rgb_reg = 3'b111; end
            18'b010010011100000011: begin rgb_reg = 3'b111; end
            18'b010010011100000100: begin rgb_reg = 3'b111; end
            18'b010010011100000101: begin rgb_reg = 3'b111; end
            18'b010010011100000110: begin rgb_reg = 3'b111; end
            18'b010010011100000111: begin rgb_reg = 3'b111; end
            18'b010010011100001000: begin rgb_reg = 3'b111; end
            18'b010010011100001001: begin rgb_reg = 3'b111; end
            18'b010010011100001010: begin rgb_reg = 3'b111; end
            18'b010010011100001011: begin rgb_reg = 3'b111; end
            18'b010010011100001100: begin rgb_reg = 3'b111; end
            18'b010010011100010011: begin rgb_reg = 3'b111; end
            18'b010010011100010100: begin rgb_reg = 3'b111; end
            18'b010010011100010101: begin rgb_reg = 3'b111; end
            18'b010010011100011110: begin rgb_reg = 3'b111; end
            18'b010010011100011111: begin rgb_reg = 3'b111; end
            18'b010010011100100000: begin rgb_reg = 3'b111; end
            18'b010010011100100001: begin rgb_reg = 3'b111; end
            18'b010010011100100010: begin rgb_reg = 3'b111; end
            18'b010010011100100011: begin rgb_reg = 3'b111; end
            18'b010010011100100100: begin rgb_reg = 3'b111; end
            18'b010010011100101100: begin rgb_reg = 3'b111; end
            18'b010010011100101101: begin rgb_reg = 3'b111; end
            18'b010010011100101110: begin rgb_reg = 3'b111; end
            18'b010010011100101111: begin rgb_reg = 3'b111; end
            18'b010010011100110000: begin rgb_reg = 3'b111; end
            18'b010010011100110001: begin rgb_reg = 3'b111; end
            18'b010010011100110010: begin rgb_reg = 3'b111; end
            18'b010010011100111100: begin rgb_reg = 3'b111; end
            18'b010010011100111101: begin rgb_reg = 3'b111; end
            18'b010010100011000000: begin rgb_reg = 3'b111; end
            18'b010010100011000001: begin rgb_reg = 3'b111; end
            18'b010010100011001011: begin rgb_reg = 3'b111; end
            18'b010010100011001100: begin rgb_reg = 3'b111; end
            18'b010010100011001101: begin rgb_reg = 3'b111; end
            18'b010010100011010100: begin rgb_reg = 3'b111; end
            18'b010010100011010101: begin rgb_reg = 3'b111; end
            18'b010010100011011001: begin rgb_reg = 3'b111; end
            18'b010010100011011010: begin rgb_reg = 3'b111; end
            18'b010010100011100010: begin rgb_reg = 3'b111; end
            18'b010010100011100011: begin rgb_reg = 3'b111; end
            18'b010010100011101001: begin rgb_reg = 3'b111; end
            18'b010010100011101010: begin rgb_reg = 3'b111; end
            18'b010010100011101011: begin rgb_reg = 3'b111; end
            18'b010010100011101100: begin rgb_reg = 3'b111; end
            18'b010010100011110100: begin rgb_reg = 3'b111; end
            18'b010010100011110101: begin rgb_reg = 3'b111; end
            18'b010010100011111101: begin rgb_reg = 3'b111; end
            18'b010010100011111110: begin rgb_reg = 3'b111; end
            18'b010010100100000001: begin rgb_reg = 3'b111; end
            18'b010010100100000010: begin rgb_reg = 3'b111; end
            18'b010010100100000011: begin rgb_reg = 3'b111; end
            18'b010010100100010001: begin rgb_reg = 3'b111; end
            18'b010010100100010010: begin rgb_reg = 3'b111; end
            18'b010010100100010011: begin rgb_reg = 3'b111; end
            18'b010010100100010100: begin rgb_reg = 3'b111; end
            18'b010010100100010101: begin rgb_reg = 3'b111; end
            18'b010010100100011100: begin rgb_reg = 3'b111; end
            18'b010010100100011101: begin rgb_reg = 3'b111; end
            18'b010010100100011110: begin rgb_reg = 3'b111; end
            18'b010010100100100101: begin rgb_reg = 3'b111; end
            18'b010010100100100110: begin rgb_reg = 3'b111; end
            18'b010010100100101010: begin rgb_reg = 3'b111; end
            18'b010010100100101011: begin rgb_reg = 3'b111; end
            18'b010010100100110011: begin rgb_reg = 3'b111; end
            18'b010010100100110100: begin rgb_reg = 3'b111; end
            18'b010010100100111010: begin rgb_reg = 3'b111; end
            18'b010010100100111011: begin rgb_reg = 3'b111; end
            18'b010010100100111100: begin rgb_reg = 3'b111; end
            18'b010010100100111101: begin rgb_reg = 3'b111; end
            18'b010010101011000000: begin rgb_reg = 3'b111; end
            18'b010010101011000001: begin rgb_reg = 3'b111; end
            18'b010010101011001011: begin rgb_reg = 3'b111; end
            18'b010010101011001100: begin rgb_reg = 3'b111; end
            18'b010010101011001101: begin rgb_reg = 3'b111; end
            18'b010010101011010100: begin rgb_reg = 3'b111; end
            18'b010010101011010101: begin rgb_reg = 3'b111; end
            18'b010010101011010110: begin rgb_reg = 3'b111; end
            18'b010010101011011001: begin rgb_reg = 3'b111; end
            18'b010010101011011010: begin rgb_reg = 3'b111; end
            18'b010010101011100010: begin rgb_reg = 3'b111; end
            18'b010010101011100011: begin rgb_reg = 3'b111; end
            18'b010010101011101000: begin rgb_reg = 3'b111; end
            18'b010010101011101001: begin rgb_reg = 3'b111; end
            18'b010010101011101010: begin rgb_reg = 3'b111; end
            18'b010010101011101011: begin rgb_reg = 3'b111; end
            18'b010010101011101100: begin rgb_reg = 3'b111; end
            18'b010010101011110100: begin rgb_reg = 3'b111; end
            18'b010010101011110101: begin rgb_reg = 3'b111; end
            18'b010010101011111101: begin rgb_reg = 3'b111; end
            18'b010010101011111110: begin rgb_reg = 3'b111; end
            18'b010010101100000001: begin rgb_reg = 3'b111; end
            18'b010010101100000010: begin rgb_reg = 3'b111; end
            18'b010010101100000011: begin rgb_reg = 3'b111; end
            18'b010010101100010001: begin rgb_reg = 3'b111; end
            18'b010010101100010010: begin rgb_reg = 3'b111; end
            18'b010010101100010011: begin rgb_reg = 3'b111; end
            18'b010010101100010100: begin rgb_reg = 3'b111; end
            18'b010010101100010101: begin rgb_reg = 3'b111; end
            18'b010010101100011100: begin rgb_reg = 3'b111; end
            18'b010010101100011101: begin rgb_reg = 3'b111; end
            18'b010010101100011110: begin rgb_reg = 3'b111; end
            18'b010010101100100101: begin rgb_reg = 3'b111; end
            18'b010010101100100110: begin rgb_reg = 3'b111; end
            18'b010010101100100111: begin rgb_reg = 3'b111; end
            18'b010010101100101010: begin rgb_reg = 3'b111; end
            18'b010010101100101011: begin rgb_reg = 3'b111; end
            18'b010010101100110011: begin rgb_reg = 3'b111; end
            18'b010010101100110100: begin rgb_reg = 3'b111; end
            18'b010010101100111001: begin rgb_reg = 3'b111; end
            18'b010010101100111010: begin rgb_reg = 3'b111; end
            18'b010010101100111011: begin rgb_reg = 3'b111; end
            18'b010010101100111100: begin rgb_reg = 3'b111; end
            18'b010010101100111101: begin rgb_reg = 3'b111; end
            18'b010010110010111110: begin rgb_reg = 3'b111; end
            18'b010010110010111111: begin rgb_reg = 3'b111; end
            18'b010010110011000000: begin rgb_reg = 3'b111; end
            18'b010010110011000001: begin rgb_reg = 3'b111; end
            18'b010010110011001011: begin rgb_reg = 3'b111; end
            18'b010010110011001100: begin rgb_reg = 3'b111; end
            18'b010010110011001101: begin rgb_reg = 3'b111; end
            18'b010010110011010010: begin rgb_reg = 3'b111; end
            18'b010010110011010011: begin rgb_reg = 3'b111; end
            18'b010010110011010100: begin rgb_reg = 3'b111; end
            18'b010010110011010101: begin rgb_reg = 3'b111; end
            18'b010010110011010110: begin rgb_reg = 3'b111; end
            18'b010010110011011001: begin rgb_reg = 3'b111; end
            18'b010010110011011010: begin rgb_reg = 3'b111; end
            18'b010010110011100010: begin rgb_reg = 3'b111; end
            18'b010010110011100011: begin rgb_reg = 3'b111; end
            18'b010010110011101001: begin rgb_reg = 3'b111; end
            18'b010010110011101010: begin rgb_reg = 3'b111; end
            18'b010010110011101011: begin rgb_reg = 3'b111; end
            18'b010010110011101100: begin rgb_reg = 3'b111; end
            18'b010010110011110100: begin rgb_reg = 3'b111; end
            18'b010010110011110101: begin rgb_reg = 3'b111; end
            18'b010010110011111011: begin rgb_reg = 3'b111; end
            18'b010010110011111100: begin rgb_reg = 3'b111; end
            18'b010010110011111101: begin rgb_reg = 3'b111; end
            18'b010010110011111110: begin rgb_reg = 3'b111; end
            18'b010010110100000001: begin rgb_reg = 3'b111; end
            18'b010010110100000010: begin rgb_reg = 3'b111; end
            18'b010010110100000011: begin rgb_reg = 3'b111; end
            18'b010010110100000100: begin rgb_reg = 3'b111; end
            18'b010010110100000101: begin rgb_reg = 3'b111; end
            18'b010010110100000110: begin rgb_reg = 3'b111; end
            18'b010010110100000111: begin rgb_reg = 3'b111; end
            18'b010010110100001000: begin rgb_reg = 3'b111; end
            18'b010010110100001001: begin rgb_reg = 3'b111; end
            18'b010010110100010001: begin rgb_reg = 3'b111; end
            18'b010010110100010010: begin rgb_reg = 3'b111; end
            18'b010010110100010011: begin rgb_reg = 3'b111; end
            18'b010010110100010100: begin rgb_reg = 3'b111; end
            18'b010010110100010101: begin rgb_reg = 3'b111; end
            18'b010010110100011100: begin rgb_reg = 3'b111; end
            18'b010010110100011101: begin rgb_reg = 3'b111; end
            18'b010010110100011110: begin rgb_reg = 3'b111; end
            18'b010010110100100101: begin rgb_reg = 3'b111; end
            18'b010010110100100110: begin rgb_reg = 3'b111; end
            18'b010010110100100111: begin rgb_reg = 3'b111; end
            18'b010010110100101010: begin rgb_reg = 3'b111; end
            18'b010010110100101011: begin rgb_reg = 3'b111; end
            18'b010010110100110011: begin rgb_reg = 3'b111; end
            18'b010010110100110100: begin rgb_reg = 3'b111; end
            18'b010010110100111010: begin rgb_reg = 3'b111; end
            18'b010010110100111011: begin rgb_reg = 3'b111; end
            18'b010010110100111100: begin rgb_reg = 3'b111; end
            18'b010010110100111101: begin rgb_reg = 3'b111; end
            18'b010010111010111110: begin rgb_reg = 3'b111; end
            18'b010010111010111111: begin rgb_reg = 3'b111; end
            18'b010010111011001011: begin rgb_reg = 3'b111; end
            18'b010010111011001100: begin rgb_reg = 3'b111; end
            18'b010010111011001101: begin rgb_reg = 3'b111; end
            18'b010010111011010010: begin rgb_reg = 3'b111; end
            18'b010010111011010011: begin rgb_reg = 3'b111; end
            18'b010010111011010100: begin rgb_reg = 3'b111; end
            18'b010010111011010101: begin rgb_reg = 3'b111; end
            18'b010010111011010110: begin rgb_reg = 3'b111; end
            18'b010010111011100010: begin rgb_reg = 3'b111; end
            18'b010010111011100011: begin rgb_reg = 3'b111; end
            18'b010010111011101011: begin rgb_reg = 3'b111; end
            18'b010010111011101100: begin rgb_reg = 3'b111; end
            18'b010010111011110100: begin rgb_reg = 3'b111; end
            18'b010010111011110101: begin rgb_reg = 3'b111; end
            18'b010010111011111010: begin rgb_reg = 3'b111; end
            18'b010010111011111011: begin rgb_reg = 3'b111; end
            18'b010010111011111100: begin rgb_reg = 3'b111; end
            18'b010010111011111101: begin rgb_reg = 3'b111; end
            18'b010010111011111110: begin rgb_reg = 3'b111; end
            18'b010010111100000001: begin rgb_reg = 3'b111; end
            18'b010010111100000010: begin rgb_reg = 3'b111; end
            18'b010010111100000011: begin rgb_reg = 3'b111; end
            18'b010010111100000100: begin rgb_reg = 3'b111; end
            18'b010010111100000101: begin rgb_reg = 3'b111; end
            18'b010010111100000110: begin rgb_reg = 3'b111; end
            18'b010010111100000111: begin rgb_reg = 3'b111; end
            18'b010010111100001000: begin rgb_reg = 3'b111; end
            18'b010010111100001001: begin rgb_reg = 3'b111; end
            18'b010010111100010011: begin rgb_reg = 3'b111; end
            18'b010010111100010100: begin rgb_reg = 3'b111; end
            18'b010010111100010101: begin rgb_reg = 3'b111; end
            18'b010010111100011100: begin rgb_reg = 3'b111; end
            18'b010010111100011101: begin rgb_reg = 3'b111; end
            18'b010010111100011110: begin rgb_reg = 3'b111; end
            18'b010010111100100101: begin rgb_reg = 3'b111; end
            18'b010010111100100110: begin rgb_reg = 3'b111; end
            18'b010010111100100111: begin rgb_reg = 3'b111; end
            18'b010010111100110011: begin rgb_reg = 3'b111; end
            18'b010010111100110100: begin rgb_reg = 3'b111; end
            18'b010010111100111100: begin rgb_reg = 3'b111; end
            18'b010010111100111101: begin rgb_reg = 3'b111; end
            18'b010011000010111110: begin rgb_reg = 3'b111; end
            18'b010011000010111111: begin rgb_reg = 3'b111; end
            18'b010011000011001011: begin rgb_reg = 3'b111; end
            18'b010011000011001100: begin rgb_reg = 3'b111; end
            18'b010011000011001101: begin rgb_reg = 3'b111; end
            18'b010011000011010010: begin rgb_reg = 3'b111; end
            18'b010011000011010011: begin rgb_reg = 3'b111; end
            18'b010011000011010100: begin rgb_reg = 3'b111; end
            18'b010011000011010101: begin rgb_reg = 3'b111; end
            18'b010011000011010110: begin rgb_reg = 3'b111; end
            18'b010011000011100010: begin rgb_reg = 3'b111; end
            18'b010011000011100011: begin rgb_reg = 3'b111; end
            18'b010011000011101011: begin rgb_reg = 3'b111; end
            18'b010011000011101100: begin rgb_reg = 3'b111; end
            18'b010011000011110100: begin rgb_reg = 3'b111; end
            18'b010011000011110101: begin rgb_reg = 3'b111; end
            18'b010011000011111010: begin rgb_reg = 3'b111; end
            18'b010011000011111011: begin rgb_reg = 3'b111; end
            18'b010011000011111100: begin rgb_reg = 3'b111; end
            18'b010011000011111101: begin rgb_reg = 3'b111; end
            18'b010011000011111110: begin rgb_reg = 3'b111; end
            18'b010011000100000001: begin rgb_reg = 3'b111; end
            18'b010011000100000010: begin rgb_reg = 3'b111; end
            18'b010011000100000011: begin rgb_reg = 3'b111; end
            18'b010011000100000100: begin rgb_reg = 3'b111; end
            18'b010011000100000101: begin rgb_reg = 3'b111; end
            18'b010011000100000110: begin rgb_reg = 3'b111; end
            18'b010011000100000111: begin rgb_reg = 3'b111; end
            18'b010011000100001000: begin rgb_reg = 3'b111; end
            18'b010011000100001001: begin rgb_reg = 3'b111; end
            18'b010011000100010011: begin rgb_reg = 3'b111; end
            18'b010011000100010100: begin rgb_reg = 3'b111; end
            18'b010011000100010101: begin rgb_reg = 3'b111; end
            18'b010011000100011100: begin rgb_reg = 3'b111; end
            18'b010011000100011101: begin rgb_reg = 3'b111; end
            18'b010011000100011110: begin rgb_reg = 3'b111; end
            18'b010011000100100101: begin rgb_reg = 3'b111; end
            18'b010011000100100110: begin rgb_reg = 3'b111; end
            18'b010011000100110011: begin rgb_reg = 3'b111; end
            18'b010011000100110100: begin rgb_reg = 3'b111; end
            18'b010011000100111100: begin rgb_reg = 3'b111; end
            18'b010011000100111101: begin rgb_reg = 3'b111; end
            18'b010011001010111110: begin rgb_reg = 3'b111; end
            18'b010011001010111111: begin rgb_reg = 3'b111; end
            18'b010011001011000000: begin rgb_reg = 3'b111; end
            18'b010011001011000001: begin rgb_reg = 3'b111; end
            18'b010011001011000010: begin rgb_reg = 3'b111; end
            18'b010011001011000011: begin rgb_reg = 3'b111; end
            18'b010011001011000100: begin rgb_reg = 3'b111; end
            18'b010011001011000101: begin rgb_reg = 3'b111; end
            18'b010011001011000110: begin rgb_reg = 3'b111; end
            18'b010011001011001011: begin rgb_reg = 3'b111; end
            18'b010011001011001100: begin rgb_reg = 3'b111; end
            18'b010011001011001101: begin rgb_reg = 3'b111; end
            18'b010011001011010000: begin rgb_reg = 3'b111; end
            18'b010011001011010001: begin rgb_reg = 3'b111; end
            18'b010011001011010100: begin rgb_reg = 3'b111; end
            18'b010011001011010101: begin rgb_reg = 3'b111; end
            18'b010011001011010110: begin rgb_reg = 3'b111; end
            18'b010011001011011101: begin rgb_reg = 3'b111; end
            18'b010011001011011110: begin rgb_reg = 3'b111; end
            18'b010011001011011111: begin rgb_reg = 3'b111; end
            18'b010011001011100000: begin rgb_reg = 3'b111; end
            18'b010011001011100001: begin rgb_reg = 3'b111; end
            18'b010011001011101011: begin rgb_reg = 3'b111; end
            18'b010011001011101100: begin rgb_reg = 3'b111; end
            18'b010011001011110100: begin rgb_reg = 3'b111; end
            18'b010011001011110101: begin rgb_reg = 3'b111; end
            18'b010011001011111000: begin rgb_reg = 3'b111; end
            18'b010011001011111001: begin rgb_reg = 3'b111; end
            18'b010011001011111010: begin rgb_reg = 3'b111; end
            18'b010011001011111101: begin rgb_reg = 3'b111; end
            18'b010011001011111110: begin rgb_reg = 3'b111; end
            18'b010011001100001010: begin rgb_reg = 3'b111; end
            18'b010011001100001011: begin rgb_reg = 3'b111; end
            18'b010011001100001100: begin rgb_reg = 3'b111; end
            18'b010011001100010011: begin rgb_reg = 3'b111; end
            18'b010011001100010100: begin rgb_reg = 3'b111; end
            18'b010011001100010101: begin rgb_reg = 3'b111; end
            18'b010011001100011110: begin rgb_reg = 3'b111; end
            18'b010011001100011111: begin rgb_reg = 3'b111; end
            18'b010011001100100000: begin rgb_reg = 3'b111; end
            18'b010011001100100001: begin rgb_reg = 3'b111; end
            18'b010011001100100010: begin rgb_reg = 3'b111; end
            18'b010011001100100011: begin rgb_reg = 3'b111; end
            18'b010011001100100100: begin rgb_reg = 3'b111; end
            18'b010011001100101110: begin rgb_reg = 3'b111; end
            18'b010011001100101111: begin rgb_reg = 3'b111; end
            18'b010011001100110000: begin rgb_reg = 3'b111; end
            18'b010011001100110001: begin rgb_reg = 3'b111; end
            18'b010011001100110010: begin rgb_reg = 3'b111; end
            18'b010011001100111100: begin rgb_reg = 3'b111; end
            18'b010011001100111101: begin rgb_reg = 3'b111; end
            18'b010011010010111110: begin rgb_reg = 3'b111; end
            18'b010011010010111111: begin rgb_reg = 3'b111; end
            18'b010011010011000000: begin rgb_reg = 3'b111; end
            18'b010011010011000001: begin rgb_reg = 3'b111; end
            18'b010011010011000010: begin rgb_reg = 3'b111; end
            18'b010011010011000011: begin rgb_reg = 3'b111; end
            18'b010011010011000100: begin rgb_reg = 3'b111; end
            18'b010011010011000101: begin rgb_reg = 3'b111; end
            18'b010011010011000110: begin rgb_reg = 3'b111; end
            18'b010011010011001011: begin rgb_reg = 3'b111; end
            18'b010011010011001100: begin rgb_reg = 3'b111; end
            18'b010011010011001101: begin rgb_reg = 3'b111; end
            18'b010011010011010000: begin rgb_reg = 3'b111; end
            18'b010011010011010001: begin rgb_reg = 3'b111; end
            18'b010011010011010100: begin rgb_reg = 3'b111; end
            18'b010011010011010101: begin rgb_reg = 3'b111; end
            18'b010011010011010110: begin rgb_reg = 3'b111; end
            18'b010011010011011101: begin rgb_reg = 3'b111; end
            18'b010011010011011110: begin rgb_reg = 3'b111; end
            18'b010011010011011111: begin rgb_reg = 3'b111; end
            18'b010011010011100000: begin rgb_reg = 3'b111; end
            18'b010011010011100001: begin rgb_reg = 3'b111; end
            18'b010011010011101011: begin rgb_reg = 3'b111; end
            18'b010011010011101100: begin rgb_reg = 3'b111; end
            18'b010011010011110100: begin rgb_reg = 3'b111; end
            18'b010011010011110101: begin rgb_reg = 3'b111; end
            18'b010011010011111000: begin rgb_reg = 3'b111; end
            18'b010011010011111001: begin rgb_reg = 3'b111; end
            18'b010011010011111010: begin rgb_reg = 3'b111; end
            18'b010011010011111101: begin rgb_reg = 3'b111; end
            18'b010011010011111110: begin rgb_reg = 3'b111; end
            18'b010011010100001010: begin rgb_reg = 3'b111; end
            18'b010011010100001011: begin rgb_reg = 3'b111; end
            18'b010011010100001100: begin rgb_reg = 3'b111; end
            18'b010011010100010011: begin rgb_reg = 3'b111; end
            18'b010011010100010100: begin rgb_reg = 3'b111; end
            18'b010011010100010101: begin rgb_reg = 3'b111; end
            18'b010011010100011110: begin rgb_reg = 3'b111; end
            18'b010011010100011111: begin rgb_reg = 3'b111; end
            18'b010011010100100000: begin rgb_reg = 3'b111; end
            18'b010011010100100001: begin rgb_reg = 3'b111; end
            18'b010011010100100010: begin rgb_reg = 3'b111; end
            18'b010011010100100011: begin rgb_reg = 3'b111; end
            18'b010011010100100100: begin rgb_reg = 3'b111; end
            18'b010011010100101110: begin rgb_reg = 3'b111; end
            18'b010011010100101111: begin rgb_reg = 3'b111; end
            18'b010011010100110000: begin rgb_reg = 3'b111; end
            18'b010011010100110001: begin rgb_reg = 3'b111; end
            18'b010011010100110010: begin rgb_reg = 3'b111; end
            18'b010011010100111100: begin rgb_reg = 3'b111; end
            18'b010011010100111101: begin rgb_reg = 3'b111; end
            18'b010011011010111110: begin rgb_reg = 3'b111; end
            18'b010011011010111111: begin rgb_reg = 3'b111; end
            18'b010011011011000111: begin rgb_reg = 3'b111; end
            18'b010011011011001000: begin rgb_reg = 3'b111; end
            18'b010011011011001011: begin rgb_reg = 3'b111; end
            18'b010011011011001100: begin rgb_reg = 3'b111; end
            18'b010011011011001101: begin rgb_reg = 3'b111; end
            18'b010011011011001110: begin rgb_reg = 3'b111; end
            18'b010011011011001111: begin rgb_reg = 3'b111; end
            18'b010011011011010100: begin rgb_reg = 3'b111; end
            18'b010011011011010101: begin rgb_reg = 3'b111; end
            18'b010011011011010110: begin rgb_reg = 3'b111; end
            18'b010011011011100010: begin rgb_reg = 3'b111; end
            18'b010011011011100011: begin rgb_reg = 3'b111; end
            18'b010011011011101011: begin rgb_reg = 3'b111; end
            18'b010011011011101100: begin rgb_reg = 3'b111; end
            18'b010011011011110100: begin rgb_reg = 3'b111; end
            18'b010011011011110101: begin rgb_reg = 3'b111; end
            18'b010011011011110110: begin rgb_reg = 3'b111; end
            18'b010011011011110111: begin rgb_reg = 3'b111; end
            18'b010011011011111101: begin rgb_reg = 3'b111; end
            18'b010011011011111110: begin rgb_reg = 3'b111; end
            18'b010011011100001010: begin rgb_reg = 3'b111; end
            18'b010011011100001011: begin rgb_reg = 3'b111; end
            18'b010011011100001100: begin rgb_reg = 3'b111; end
            18'b010011011100010011: begin rgb_reg = 3'b111; end
            18'b010011011100010100: begin rgb_reg = 3'b111; end
            18'b010011011100010101: begin rgb_reg = 3'b111; end
            18'b010011011100011100: begin rgb_reg = 3'b111; end
            18'b010011011100011101: begin rgb_reg = 3'b111; end
            18'b010011011100011110: begin rgb_reg = 3'b111; end
            18'b010011011100100101: begin rgb_reg = 3'b111; end
            18'b010011011100100110: begin rgb_reg = 3'b111; end
            18'b010011011100100111: begin rgb_reg = 3'b111; end
            18'b010011011100101100: begin rgb_reg = 3'b111; end
            18'b010011011100101101: begin rgb_reg = 3'b111; end
            18'b010011011100111100: begin rgb_reg = 3'b111; end
            18'b010011011100111101: begin rgb_reg = 3'b111; end
            18'b010011100010111110: begin rgb_reg = 3'b111; end
            18'b010011100010111111: begin rgb_reg = 3'b111; end
            18'b010011100011000111: begin rgb_reg = 3'b111; end
            18'b010011100011001000: begin rgb_reg = 3'b111; end
            18'b010011100011001011: begin rgb_reg = 3'b111; end
            18'b010011100011001100: begin rgb_reg = 3'b111; end
            18'b010011100011001101: begin rgb_reg = 3'b111; end
            18'b010011100011001110: begin rgb_reg = 3'b111; end
            18'b010011100011001111: begin rgb_reg = 3'b111; end
            18'b010011100011010100: begin rgb_reg = 3'b111; end
            18'b010011100011010101: begin rgb_reg = 3'b111; end
            18'b010011100011010110: begin rgb_reg = 3'b111; end
            18'b010011100011100010: begin rgb_reg = 3'b111; end
            18'b010011100011100011: begin rgb_reg = 3'b111; end
            18'b010011100011101011: begin rgb_reg = 3'b111; end
            18'b010011100011101100: begin rgb_reg = 3'b111; end
            18'b010011100011110100: begin rgb_reg = 3'b111; end
            18'b010011100011110101: begin rgb_reg = 3'b111; end
            18'b010011100011110110: begin rgb_reg = 3'b111; end
            18'b010011100011110111: begin rgb_reg = 3'b111; end
            18'b010011100011111101: begin rgb_reg = 3'b111; end
            18'b010011100011111110: begin rgb_reg = 3'b111; end
            18'b010011100100001010: begin rgb_reg = 3'b111; end
            18'b010011100100001011: begin rgb_reg = 3'b111; end
            18'b010011100100001100: begin rgb_reg = 3'b111; end
            18'b010011100100010011: begin rgb_reg = 3'b111; end
            18'b010011100100010100: begin rgb_reg = 3'b111; end
            18'b010011100100010101: begin rgb_reg = 3'b111; end
            18'b010011100100011100: begin rgb_reg = 3'b111; end
            18'b010011100100011101: begin rgb_reg = 3'b111; end
            18'b010011100100011110: begin rgb_reg = 3'b111; end
            18'b010011100100100101: begin rgb_reg = 3'b111; end
            18'b010011100100100110: begin rgb_reg = 3'b111; end
            18'b010011100100100111: begin rgb_reg = 3'b111; end
            18'b010011100100101100: begin rgb_reg = 3'b111; end
            18'b010011100100101101: begin rgb_reg = 3'b111; end
            18'b010011100100111100: begin rgb_reg = 3'b111; end
            18'b010011100100111101: begin rgb_reg = 3'b111; end
            18'b010011101010111110: begin rgb_reg = 3'b111; end
            18'b010011101010111111: begin rgb_reg = 3'b111; end
            18'b010011101011000111: begin rgb_reg = 3'b111; end
            18'b010011101011001000: begin rgb_reg = 3'b111; end
            18'b010011101011001011: begin rgb_reg = 3'b111; end
            18'b010011101011001100: begin rgb_reg = 3'b111; end
            18'b010011101011001101: begin rgb_reg = 3'b111; end
            18'b010011101011010100: begin rgb_reg = 3'b111; end
            18'b010011101011010101: begin rgb_reg = 3'b111; end
            18'b010011101011010110: begin rgb_reg = 3'b111; end
            18'b010011101011011001: begin rgb_reg = 3'b111; end
            18'b010011101011011010: begin rgb_reg = 3'b111; end
            18'b010011101011100010: begin rgb_reg = 3'b111; end
            18'b010011101011100011: begin rgb_reg = 3'b111; end
            18'b010011101011101011: begin rgb_reg = 3'b111; end
            18'b010011101011101100: begin rgb_reg = 3'b111; end
            18'b010011101011110100: begin rgb_reg = 3'b111; end
            18'b010011101011110101: begin rgb_reg = 3'b111; end
            18'b010011101011111101: begin rgb_reg = 3'b111; end
            18'b010011101011111110: begin rgb_reg = 3'b111; end
            18'b010011101100000001: begin rgb_reg = 3'b111; end
            18'b010011101100000010: begin rgb_reg = 3'b111; end
            18'b010011101100001010: begin rgb_reg = 3'b111; end
            18'b010011101100001011: begin rgb_reg = 3'b111; end
            18'b010011101100001100: begin rgb_reg = 3'b111; end
            18'b010011101100010011: begin rgb_reg = 3'b111; end
            18'b010011101100010100: begin rgb_reg = 3'b111; end
            18'b010011101100010101: begin rgb_reg = 3'b111; end
            18'b010011101100011100: begin rgb_reg = 3'b111; end
            18'b010011101100011101: begin rgb_reg = 3'b111; end
            18'b010011101100011110: begin rgb_reg = 3'b111; end
            18'b010011101100100101: begin rgb_reg = 3'b111; end
            18'b010011101100100110: begin rgb_reg = 3'b111; end
            18'b010011101100100111: begin rgb_reg = 3'b111; end
            18'b010011101100101010: begin rgb_reg = 3'b111; end
            18'b010011101100101011: begin rgb_reg = 3'b111; end
            18'b010011101100111100: begin rgb_reg = 3'b111; end
            18'b010011101100111101: begin rgb_reg = 3'b111; end
            18'b010011110010111110: begin rgb_reg = 3'b111; end
            18'b010011110010111111: begin rgb_reg = 3'b111; end
            18'b010011110011000111: begin rgb_reg = 3'b111; end
            18'b010011110011001000: begin rgb_reg = 3'b111; end
            18'b010011110011001011: begin rgb_reg = 3'b111; end
            18'b010011110011001100: begin rgb_reg = 3'b111; end
            18'b010011110011001101: begin rgb_reg = 3'b111; end
            18'b010011110011010100: begin rgb_reg = 3'b111; end
            18'b010011110011010101: begin rgb_reg = 3'b111; end
            18'b010011110011010110: begin rgb_reg = 3'b111; end
            18'b010011110011011001: begin rgb_reg = 3'b111; end
            18'b010011110011011010: begin rgb_reg = 3'b111; end
            18'b010011110011100010: begin rgb_reg = 3'b111; end
            18'b010011110011100011: begin rgb_reg = 3'b111; end
            18'b010011110011101011: begin rgb_reg = 3'b111; end
            18'b010011110011101100: begin rgb_reg = 3'b111; end
            18'b010011110011110100: begin rgb_reg = 3'b111; end
            18'b010011110011110101: begin rgb_reg = 3'b111; end
            18'b010011110011111101: begin rgb_reg = 3'b111; end
            18'b010011110011111110: begin rgb_reg = 3'b111; end
            18'b010011110100000001: begin rgb_reg = 3'b111; end
            18'b010011110100000010: begin rgb_reg = 3'b111; end
            18'b010011110100000011: begin rgb_reg = 3'b111; end
            18'b010011110100001010: begin rgb_reg = 3'b111; end
            18'b010011110100001011: begin rgb_reg = 3'b111; end
            18'b010011110100001100: begin rgb_reg = 3'b111; end
            18'b010011110100010011: begin rgb_reg = 3'b111; end
            18'b010011110100010100: begin rgb_reg = 3'b111; end
            18'b010011110100010101: begin rgb_reg = 3'b111; end
            18'b010011110100011100: begin rgb_reg = 3'b111; end
            18'b010011110100011101: begin rgb_reg = 3'b111; end
            18'b010011110100011110: begin rgb_reg = 3'b111; end
            18'b010011110100100101: begin rgb_reg = 3'b111; end
            18'b010011110100100110: begin rgb_reg = 3'b111; end
            18'b010011110100100111: begin rgb_reg = 3'b111; end
            18'b010011110100101010: begin rgb_reg = 3'b111; end
            18'b010011110100101011: begin rgb_reg = 3'b111; end
            18'b010011110100111100: begin rgb_reg = 3'b111; end
            18'b010011110100111101: begin rgb_reg = 3'b111; end
            18'b010011111010111110: begin rgb_reg = 3'b111; end
            18'b010011111010111111: begin rgb_reg = 3'b111; end
            18'b010011111011000000: begin rgb_reg = 3'b111; end
            18'b010011111011000001: begin rgb_reg = 3'b111; end
            18'b010011111011000010: begin rgb_reg = 3'b111; end
            18'b010011111011000011: begin rgb_reg = 3'b111; end
            18'b010011111011000100: begin rgb_reg = 3'b111; end
            18'b010011111011000101: begin rgb_reg = 3'b111; end
            18'b010011111011000110: begin rgb_reg = 3'b111; end
            18'b010011111011000111: begin rgb_reg = 3'b111; end
            18'b010011111011001000: begin rgb_reg = 3'b111; end
            18'b010011111011001100: begin rgb_reg = 3'b111; end
            18'b010011111011001101: begin rgb_reg = 3'b111; end
            18'b010011111011001110: begin rgb_reg = 3'b111; end
            18'b010011111011001111: begin rgb_reg = 3'b111; end
            18'b010011111011010000: begin rgb_reg = 3'b111; end
            18'b010011111011010001: begin rgb_reg = 3'b111; end
            18'b010011111011010010: begin rgb_reg = 3'b111; end
            18'b010011111011010011: begin rgb_reg = 3'b111; end
            18'b010011111011010100: begin rgb_reg = 3'b111; end
            18'b010011111011010101: begin rgb_reg = 3'b111; end
            18'b010011111011011001: begin rgb_reg = 3'b111; end
            18'b010011111011011010: begin rgb_reg = 3'b111; end
            18'b010011111011011011: begin rgb_reg = 3'b111; end
            18'b010011111011011100: begin rgb_reg = 3'b111; end
            18'b010011111011011101: begin rgb_reg = 3'b111; end
            18'b010011111011011110: begin rgb_reg = 3'b111; end
            18'b010011111011011111: begin rgb_reg = 3'b111; end
            18'b010011111011100000: begin rgb_reg = 3'b111; end
            18'b010011111011100001: begin rgb_reg = 3'b111; end
            18'b010011111011100010: begin rgb_reg = 3'b111; end
            18'b010011111011100011: begin rgb_reg = 3'b111; end
            18'b010011111011100111: begin rgb_reg = 3'b111; end
            18'b010011111011101000: begin rgb_reg = 3'b111; end
            18'b010011111011101001: begin rgb_reg = 3'b111; end
            18'b010011111011101010: begin rgb_reg = 3'b111; end
            18'b010011111011101011: begin rgb_reg = 3'b111; end
            18'b010011111011101100: begin rgb_reg = 3'b111; end
            18'b010011111011101101: begin rgb_reg = 3'b111; end
            18'b010011111011101110: begin rgb_reg = 3'b111; end
            18'b010011111011101111: begin rgb_reg = 3'b111; end
            18'b010011111011110000: begin rgb_reg = 3'b111; end
            18'b010011111011110100: begin rgb_reg = 3'b111; end
            18'b010011111011110101: begin rgb_reg = 3'b111; end
            18'b010011111011110110: begin rgb_reg = 3'b111; end
            18'b010011111011110111: begin rgb_reg = 3'b111; end
            18'b010011111011111000: begin rgb_reg = 3'b111; end
            18'b010011111011111001: begin rgb_reg = 3'b111; end
            18'b010011111011111010: begin rgb_reg = 3'b111; end
            18'b010011111011111011: begin rgb_reg = 3'b111; end
            18'b010011111011111100: begin rgb_reg = 3'b111; end
            18'b010011111011111101: begin rgb_reg = 3'b111; end
            18'b010011111011111110: begin rgb_reg = 3'b111; end
            18'b010011111100000010: begin rgb_reg = 3'b111; end
            18'b010011111100000011: begin rgb_reg = 3'b111; end
            18'b010011111100000100: begin rgb_reg = 3'b111; end
            18'b010011111100000101: begin rgb_reg = 3'b111; end
            18'b010011111100000110: begin rgb_reg = 3'b111; end
            18'b010011111100000111: begin rgb_reg = 3'b111; end
            18'b010011111100001000: begin rgb_reg = 3'b111; end
            18'b010011111100001001: begin rgb_reg = 3'b111; end
            18'b010011111100001010: begin rgb_reg = 3'b111; end
            18'b010011111100001011: begin rgb_reg = 3'b111; end
            18'b010011111100001111: begin rgb_reg = 3'b111; end
            18'b010011111100010000: begin rgb_reg = 3'b111; end
            18'b010011111100010001: begin rgb_reg = 3'b111; end
            18'b010011111100010010: begin rgb_reg = 3'b111; end
            18'b010011111100010011: begin rgb_reg = 3'b111; end
            18'b010011111100010100: begin rgb_reg = 3'b111; end
            18'b010011111100010101: begin rgb_reg = 3'b111; end
            18'b010011111100010110: begin rgb_reg = 3'b111; end
            18'b010011111100010111: begin rgb_reg = 3'b111; end
            18'b010011111100011000: begin rgb_reg = 3'b111; end
            18'b010011111100011001: begin rgb_reg = 3'b111; end
            18'b010011111100011101: begin rgb_reg = 3'b111; end
            18'b010011111100011110: begin rgb_reg = 3'b111; end
            18'b010011111100011111: begin rgb_reg = 3'b111; end
            18'b010011111100100000: begin rgb_reg = 3'b111; end
            18'b010011111100100001: begin rgb_reg = 3'b111; end
            18'b010011111100100010: begin rgb_reg = 3'b111; end
            18'b010011111100100011: begin rgb_reg = 3'b111; end
            18'b010011111100100100: begin rgb_reg = 3'b111; end
            18'b010011111100100101: begin rgb_reg = 3'b111; end
            18'b010011111100100110: begin rgb_reg = 3'b111; end
            18'b010011111100101010: begin rgb_reg = 3'b111; end
            18'b010011111100101011: begin rgb_reg = 3'b111; end
            18'b010011111100101100: begin rgb_reg = 3'b111; end
            18'b010011111100101101: begin rgb_reg = 3'b111; end
            18'b010011111100101110: begin rgb_reg = 3'b111; end
            18'b010011111100101111: begin rgb_reg = 3'b111; end
            18'b010011111100110000: begin rgb_reg = 3'b111; end
            18'b010011111100110001: begin rgb_reg = 3'b111; end
            18'b010011111100110010: begin rgb_reg = 3'b111; end
            18'b010011111100110011: begin rgb_reg = 3'b111; end
            18'b010011111100110100: begin rgb_reg = 3'b111; end
            18'b010011111100111000: begin rgb_reg = 3'b111; end
            18'b010011111100111001: begin rgb_reg = 3'b111; end
            18'b010011111100111010: begin rgb_reg = 3'b111; end
            18'b010011111100111011: begin rgb_reg = 3'b111; end
            18'b010011111100111100: begin rgb_reg = 3'b111; end
            18'b010011111100111101: begin rgb_reg = 3'b111; end
            18'b010011111100111110: begin rgb_reg = 3'b111; end
            18'b010011111100111111: begin rgb_reg = 3'b111; end
            18'b010011111101000000: begin rgb_reg = 3'b111; end
            18'b010011111101000001: begin rgb_reg = 3'b111; end
            18'b010100000011000000: begin rgb_reg = 3'b111; end
            18'b010100000011000001: begin rgb_reg = 3'b111; end
            18'b010100000011000010: begin rgb_reg = 3'b111; end
            18'b010100000011000011: begin rgb_reg = 3'b111; end
            18'b010100000011000100: begin rgb_reg = 3'b111; end
            18'b010100000011000101: begin rgb_reg = 3'b111; end
            18'b010100000011000110: begin rgb_reg = 3'b111; end
            18'b010100000011001101: begin rgb_reg = 3'b111; end
            18'b010100000011001110: begin rgb_reg = 3'b111; end
            18'b010100000011001111: begin rgb_reg = 3'b111; end
            18'b010100000011010000: begin rgb_reg = 3'b111; end
            18'b010100000011010001: begin rgb_reg = 3'b111; end
            18'b010100000011010010: begin rgb_reg = 3'b111; end
            18'b010100000011010011: begin rgb_reg = 3'b111; end
            18'b010100000011011011: begin rgb_reg = 3'b111; end
            18'b010100000011011100: begin rgb_reg = 3'b111; end
            18'b010100000011011101: begin rgb_reg = 3'b111; end
            18'b010100000011011110: begin rgb_reg = 3'b111; end
            18'b010100000011011111: begin rgb_reg = 3'b111; end
            18'b010100000011100000: begin rgb_reg = 3'b111; end
            18'b010100000011100001: begin rgb_reg = 3'b111; end
            18'b010100000011100110: begin rgb_reg = 3'b111; end
            18'b010100000011100111: begin rgb_reg = 3'b111; end
            18'b010100000011101000: begin rgb_reg = 3'b111; end
            18'b010100000011101001: begin rgb_reg = 3'b111; end
            18'b010100000011101010: begin rgb_reg = 3'b111; end
            18'b010100000011101011: begin rgb_reg = 3'b111; end
            18'b010100000011101100: begin rgb_reg = 3'b111; end
            18'b010100000011101101: begin rgb_reg = 3'b111; end
            18'b010100000011101110: begin rgb_reg = 3'b111; end
            18'b010100000011101111: begin rgb_reg = 3'b111; end
            18'b010100000011110000: begin rgb_reg = 3'b111; end
            18'b010100000011110001: begin rgb_reg = 3'b111; end
            18'b010100000011110110: begin rgb_reg = 3'b111; end
            18'b010100000011110111: begin rgb_reg = 3'b111; end
            18'b010100000011111000: begin rgb_reg = 3'b111; end
            18'b010100000011111001: begin rgb_reg = 3'b111; end
            18'b010100000011111010: begin rgb_reg = 3'b111; end
            18'b010100000011111011: begin rgb_reg = 3'b111; end
            18'b010100000011111100: begin rgb_reg = 3'b111; end
            18'b010100000100000011: begin rgb_reg = 3'b111; end
            18'b010100000100000100: begin rgb_reg = 3'b111; end
            18'b010100000100000101: begin rgb_reg = 3'b111; end
            18'b010100000100000110: begin rgb_reg = 3'b111; end
            18'b010100000100000111: begin rgb_reg = 3'b111; end
            18'b010100000100001000: begin rgb_reg = 3'b111; end
            18'b010100000100001001: begin rgb_reg = 3'b111; end
            18'b010100000100001111: begin rgb_reg = 3'b111; end
            18'b010100000100010000: begin rgb_reg = 3'b111; end
            18'b010100000100010001: begin rgb_reg = 3'b111; end
            18'b010100000100010010: begin rgb_reg = 3'b111; end
            18'b010100000100010011: begin rgb_reg = 3'b111; end
            18'b010100000100010100: begin rgb_reg = 3'b111; end
            18'b010100000100010101: begin rgb_reg = 3'b111; end
            18'b010100000100010110: begin rgb_reg = 3'b111; end
            18'b010100000100010111: begin rgb_reg = 3'b111; end
            18'b010100000100011000: begin rgb_reg = 3'b111; end
            18'b010100000100011001: begin rgb_reg = 3'b111; end
            18'b010100000100011110: begin rgb_reg = 3'b111; end
            18'b010100000100011111: begin rgb_reg = 3'b111; end
            18'b010100000100100000: begin rgb_reg = 3'b111; end
            18'b010100000100100001: begin rgb_reg = 3'b111; end
            18'b010100000100100010: begin rgb_reg = 3'b111; end
            18'b010100000100100011: begin rgb_reg = 3'b111; end
            18'b010100000100100100: begin rgb_reg = 3'b111; end
            18'b010100000100101010: begin rgb_reg = 3'b111; end
            18'b010100000100101011: begin rgb_reg = 3'b111; end
            18'b010100000100101100: begin rgb_reg = 3'b111; end
            18'b010100000100101101: begin rgb_reg = 3'b111; end
            18'b010100000100101110: begin rgb_reg = 3'b111; end
            18'b010100000100101111: begin rgb_reg = 3'b111; end
            18'b010100000100110000: begin rgb_reg = 3'b111; end
            18'b010100000100110001: begin rgb_reg = 3'b111; end
            18'b010100000100110010: begin rgb_reg = 3'b111; end
            18'b010100000100110011: begin rgb_reg = 3'b111; end
            18'b010100000100110100: begin rgb_reg = 3'b111; end
            18'b010100000100110111: begin rgb_reg = 3'b111; end
            18'b010100000100111000: begin rgb_reg = 3'b111; end
            18'b010100000100111001: begin rgb_reg = 3'b111; end
            18'b010100000100111010: begin rgb_reg = 3'b111; end
            18'b010100000100111011: begin rgb_reg = 3'b111; end
            18'b010100000100111100: begin rgb_reg = 3'b111; end
            18'b010100000100111101: begin rgb_reg = 3'b111; end
            18'b010100000100111110: begin rgb_reg = 3'b111; end
            18'b010100000100111111: begin rgb_reg = 3'b111; end
            18'b010100000101000000: begin rgb_reg = 3'b111; end
            18'b010100000101000001: begin rgb_reg = 3'b111; end
            18'b010100000101000010: begin rgb_reg = 3'b111; end
            18'b010100001011000000: begin rgb_reg = 3'b111; end
            18'b010100001011000001: begin rgb_reg = 3'b111; end
            18'b010100001011000010: begin rgb_reg = 3'b111; end
            18'b010100001011000011: begin rgb_reg = 3'b111; end
            18'b010100001011000100: begin rgb_reg = 3'b111; end
            18'b010100001011000101: begin rgb_reg = 3'b111; end
            18'b010100001011000110: begin rgb_reg = 3'b111; end
            18'b010100001011001110: begin rgb_reg = 3'b111; end
            18'b010100001011001111: begin rgb_reg = 3'b111; end
            18'b010100001011010000: begin rgb_reg = 3'b111; end
            18'b010100001011010001: begin rgb_reg = 3'b111; end
            18'b010100001011010010: begin rgb_reg = 3'b111; end
            18'b010100001011010011: begin rgb_reg = 3'b111; end
            18'b010100001011011011: begin rgb_reg = 3'b111; end
            18'b010100001011011100: begin rgb_reg = 3'b111; end
            18'b010100001011011101: begin rgb_reg = 3'b111; end
            18'b010100001011011110: begin rgb_reg = 3'b111; end
            18'b010100001011011111: begin rgb_reg = 3'b111; end
            18'b010100001011100000: begin rgb_reg = 3'b111; end
            18'b010100001011100001: begin rgb_reg = 3'b111; end
            18'b010100001011100110: begin rgb_reg = 3'b111; end
            18'b010100001011100111: begin rgb_reg = 3'b111; end
            18'b010100001011101000: begin rgb_reg = 3'b111; end
            18'b010100001011101001: begin rgb_reg = 3'b111; end
            18'b010100001011101010: begin rgb_reg = 3'b111; end
            18'b010100001011101011: begin rgb_reg = 3'b111; end
            18'b010100001011101100: begin rgb_reg = 3'b111; end
            18'b010100001011101101: begin rgb_reg = 3'b111; end
            18'b010100001011101110: begin rgb_reg = 3'b111; end
            18'b010100001011101111: begin rgb_reg = 3'b111; end
            18'b010100001011110000: begin rgb_reg = 3'b111; end
            18'b010100001011110110: begin rgb_reg = 3'b111; end
            18'b010100001011110111: begin rgb_reg = 3'b111; end
            18'b010100001011111000: begin rgb_reg = 3'b111; end
            18'b010100001011111001: begin rgb_reg = 3'b111; end
            18'b010100001011111010: begin rgb_reg = 3'b111; end
            18'b010100001011111011: begin rgb_reg = 3'b111; end
            18'b010100001011111100: begin rgb_reg = 3'b111; end
            18'b010100001100000100: begin rgb_reg = 3'b111; end
            18'b010100001100000101: begin rgb_reg = 3'b111; end
            18'b010100001100000110: begin rgb_reg = 3'b111; end
            18'b010100001100000111: begin rgb_reg = 3'b111; end
            18'b010100001100001000: begin rgb_reg = 3'b111; end
            18'b010100001100001001: begin rgb_reg = 3'b111; end
            18'b010100001100001111: begin rgb_reg = 3'b111; end
            18'b010100001100010000: begin rgb_reg = 3'b111; end
            18'b010100001100010001: begin rgb_reg = 3'b111; end
            18'b010100001100010010: begin rgb_reg = 3'b111; end
            18'b010100001100010011: begin rgb_reg = 3'b111; end
            18'b010100001100010100: begin rgb_reg = 3'b111; end
            18'b010100001100010101: begin rgb_reg = 3'b111; end
            18'b010100001100010110: begin rgb_reg = 3'b111; end
            18'b010100001100010111: begin rgb_reg = 3'b111; end
            18'b010100001100011000: begin rgb_reg = 3'b111; end
            18'b010100001100011001: begin rgb_reg = 3'b111; end
            18'b010100001100011111: begin rgb_reg = 3'b111; end
            18'b010100001100100000: begin rgb_reg = 3'b111; end
            18'b010100001100100001: begin rgb_reg = 3'b111; end
            18'b010100001100100010: begin rgb_reg = 3'b111; end
            18'b010100001100100011: begin rgb_reg = 3'b111; end
            18'b010100001100100100: begin rgb_reg = 3'b111; end
            18'b010100001100101010: begin rgb_reg = 3'b111; end
            18'b010100001100101011: begin rgb_reg = 3'b111; end
            18'b010100001100101100: begin rgb_reg = 3'b111; end
            18'b010100001100101101: begin rgb_reg = 3'b111; end
            18'b010100001100101110: begin rgb_reg = 3'b111; end
            18'b010100001100101111: begin rgb_reg = 3'b111; end
            18'b010100001100110000: begin rgb_reg = 3'b111; end
            18'b010100001100110001: begin rgb_reg = 3'b111; end
            18'b010100001100110010: begin rgb_reg = 3'b111; end
            18'b010100001100110011: begin rgb_reg = 3'b111; end
            18'b010100001100110100: begin rgb_reg = 3'b111; end
            18'b010100001100110111: begin rgb_reg = 3'b111; end
            18'b010100001100111000: begin rgb_reg = 3'b111; end
            18'b010100001100111001: begin rgb_reg = 3'b111; end
            18'b010100001100111010: begin rgb_reg = 3'b111; end
            18'b010100001100111011: begin rgb_reg = 3'b111; end
            18'b010100001100111100: begin rgb_reg = 3'b111; end
            18'b010100001100111101: begin rgb_reg = 3'b111; end
            18'b010100001100111110: begin rgb_reg = 3'b111; end
            18'b010100001100111111: begin rgb_reg = 3'b111; end
            18'b010100001101000000: begin rgb_reg = 3'b111; end
            18'b010100001101000001: begin rgb_reg = 3'b111; end
            18'b010101000010110100: begin rgb_reg = 3'b111; end
            18'b010101000010110101: begin rgb_reg = 3'b111; end
            18'b010101000010111100: begin rgb_reg = 3'b111; end
            18'b010101000010111101: begin rgb_reg = 3'b111; end
            18'b010101000100001010: begin rgb_reg = 3'b111; end
            18'b010101000100001011: begin rgb_reg = 3'b111; end
            18'b010101000100011110: begin rgb_reg = 3'b111; end
            18'b010101000100011111: begin rgb_reg = 3'b111; end
            18'b010101000100100000: begin rgb_reg = 3'b111; end
            18'b010101000100100001: begin rgb_reg = 3'b111; end
            18'b010101000100100010: begin rgb_reg = 3'b111; end
            18'b010101000100100011: begin rgb_reg = 3'b111; end
            18'b010101000100100100: begin rgb_reg = 3'b111; end
            18'b010101000100100101: begin rgb_reg = 3'b111; end
            18'b010101000101000000: begin rgb_reg = 3'b111; end
            18'b010101000101000001: begin rgb_reg = 3'b111; end
            18'b010101001010110100: begin rgb_reg = 3'b111; end
            18'b010101001010110101: begin rgb_reg = 3'b111; end
            18'b010101001010111100: begin rgb_reg = 3'b111; end
            18'b010101001010111101: begin rgb_reg = 3'b111; end
            18'b010101001100001010: begin rgb_reg = 3'b111; end
            18'b010101001100001011: begin rgb_reg = 3'b111; end
            18'b010101001100011110: begin rgb_reg = 3'b111; end
            18'b010101001100011111: begin rgb_reg = 3'b111; end
            18'b010101001100100000: begin rgb_reg = 3'b111; end
            18'b010101001100100001: begin rgb_reg = 3'b111; end
            18'b010101001100100010: begin rgb_reg = 3'b111; end
            18'b010101001100100011: begin rgb_reg = 3'b111; end
            18'b010101001100100100: begin rgb_reg = 3'b111; end
            18'b010101001100100101: begin rgb_reg = 3'b111; end
            18'b010101001101000000: begin rgb_reg = 3'b111; end
            18'b010101001101000001: begin rgb_reg = 3'b111; end
            18'b010101010010110100: begin rgb_reg = 3'b111; end
            18'b010101010010110101: begin rgb_reg = 3'b111; end
            18'b010101010010111100: begin rgb_reg = 3'b111; end
            18'b010101010010111101: begin rgb_reg = 3'b111; end
            18'b010101010100001000: begin rgb_reg = 3'b111; end
            18'b010101010100001001: begin rgb_reg = 3'b111; end
            18'b010101010100001010: begin rgb_reg = 3'b111; end
            18'b010101010100001011: begin rgb_reg = 3'b111; end
            18'b010101010100001100: begin rgb_reg = 3'b111; end
            18'b010101010100001101: begin rgb_reg = 3'b111; end
            18'b010101010100011100: begin rgb_reg = 3'b111; end
            18'b010101010100011101: begin rgb_reg = 3'b111; end
            18'b010101010101000000: begin rgb_reg = 3'b111; end
            18'b010101010101000001: begin rgb_reg = 3'b111; end
            18'b010101011010110100: begin rgb_reg = 3'b111; end
            18'b010101011010110101: begin rgb_reg = 3'b111; end
            18'b010101011010111100: begin rgb_reg = 3'b111; end
            18'b010101011010111101: begin rgb_reg = 3'b111; end
            18'b010101011100001000: begin rgb_reg = 3'b111; end
            18'b010101011100001001: begin rgb_reg = 3'b111; end
            18'b010101011100001010: begin rgb_reg = 3'b111; end
            18'b010101011100001011: begin rgb_reg = 3'b111; end
            18'b010101011100001100: begin rgb_reg = 3'b111; end
            18'b010101011100001101: begin rgb_reg = 3'b111; end
            18'b010101011100011100: begin rgb_reg = 3'b111; end
            18'b010101011100011101: begin rgb_reg = 3'b111; end
            18'b010101011101000000: begin rgb_reg = 3'b111; end
            18'b010101011101000001: begin rgb_reg = 3'b111; end
            18'b010101100010110100: begin rgb_reg = 3'b111; end
            18'b010101100010110101: begin rgb_reg = 3'b111; end
            18'b010101100010111100: begin rgb_reg = 3'b111; end
            18'b010101100010111101: begin rgb_reg = 3'b111; end
            18'b010101100011000010: begin rgb_reg = 3'b111; end
            18'b010101100011000011: begin rgb_reg = 3'b111; end
            18'b010101100011000100: begin rgb_reg = 3'b111; end
            18'b010101100011000101: begin rgb_reg = 3'b111; end
            18'b010101100011000110: begin rgb_reg = 3'b111; end
            18'b010101100011000111: begin rgb_reg = 3'b111; end
            18'b010101100011001100: begin rgb_reg = 3'b111; end
            18'b010101100011001101: begin rgb_reg = 3'b111; end
            18'b010101100011010000: begin rgb_reg = 3'b111; end
            18'b010101100011010001: begin rgb_reg = 3'b111; end
            18'b010101100011010010: begin rgb_reg = 3'b111; end
            18'b010101100011010011: begin rgb_reg = 3'b111; end
            18'b010101100011011010: begin rgb_reg = 3'b111; end
            18'b010101100011011011: begin rgb_reg = 3'b111; end
            18'b010101100011011100: begin rgb_reg = 3'b111; end
            18'b010101100011011101: begin rgb_reg = 3'b111; end
            18'b010101100011011110: begin rgb_reg = 3'b111; end
            18'b010101100011011111: begin rgb_reg = 3'b111; end
            18'b010101100011100100: begin rgb_reg = 3'b111; end
            18'b010101100011100101: begin rgb_reg = 3'b111; end
            18'b010101100011101000: begin rgb_reg = 3'b111; end
            18'b010101100011101001: begin rgb_reg = 3'b111; end
            18'b010101100011101010: begin rgb_reg = 3'b111; end
            18'b010101100011101011: begin rgb_reg = 3'b111; end
            18'b010101100011110000: begin rgb_reg = 3'b111; end
            18'b010101100011110001: begin rgb_reg = 3'b111; end
            18'b010101100011110100: begin rgb_reg = 3'b111; end
            18'b010101100011110101: begin rgb_reg = 3'b111; end
            18'b010101100011110110: begin rgb_reg = 3'b111; end
            18'b010101100011110111: begin rgb_reg = 3'b111; end
            18'b010101100011111110: begin rgb_reg = 3'b111; end
            18'b010101100011111111: begin rgb_reg = 3'b111; end
            18'b010101100100000000: begin rgb_reg = 3'b111; end
            18'b010101100100000001: begin rgb_reg = 3'b111; end
            18'b010101100100000010: begin rgb_reg = 3'b111; end
            18'b010101100100000011: begin rgb_reg = 3'b111; end
            18'b010101100100001010: begin rgb_reg = 3'b111; end
            18'b010101100100001011: begin rgb_reg = 3'b111; end
            18'b010101100100011110: begin rgb_reg = 3'b111; end
            18'b010101100100011111: begin rgb_reg = 3'b111; end
            18'b010101100100100000: begin rgb_reg = 3'b111; end
            18'b010101100100100001: begin rgb_reg = 3'b111; end
            18'b010101100100100010: begin rgb_reg = 3'b111; end
            18'b010101100100100011: begin rgb_reg = 3'b111; end
            18'b010101100100101010: begin rgb_reg = 3'b111; end
            18'b010101100100101011: begin rgb_reg = 3'b111; end
            18'b010101100100101100: begin rgb_reg = 3'b111; end
            18'b010101100100101101: begin rgb_reg = 3'b111; end
            18'b010101100100101110: begin rgb_reg = 3'b111; end
            18'b010101100100101111: begin rgb_reg = 3'b111; end
            18'b010101100100110110: begin rgb_reg = 3'b111; end
            18'b010101100100110111: begin rgb_reg = 3'b111; end
            18'b010101100100111000: begin rgb_reg = 3'b111; end
            18'b010101100100111001: begin rgb_reg = 3'b111; end
            18'b010101100100111010: begin rgb_reg = 3'b111; end
            18'b010101100100111011: begin rgb_reg = 3'b111; end
            18'b010101100101000000: begin rgb_reg = 3'b111; end
            18'b010101100101000001: begin rgb_reg = 3'b111; end
            18'b010101100101001000: begin rgb_reg = 3'b111; end
            18'b010101100101001001: begin rgb_reg = 3'b111; end
            18'b010101100101001010: begin rgb_reg = 3'b111; end
            18'b010101100101001011: begin rgb_reg = 3'b111; end
            18'b010101100101001100: begin rgb_reg = 3'b111; end
            18'b010101100101001101: begin rgb_reg = 3'b111; end
            18'b010101101010110100: begin rgb_reg = 3'b111; end
            18'b010101101010110101: begin rgb_reg = 3'b111; end
            18'b010101101010111100: begin rgb_reg = 3'b111; end
            18'b010101101010111101: begin rgb_reg = 3'b111; end
            18'b010101101011000010: begin rgb_reg = 3'b111; end
            18'b010101101011000011: begin rgb_reg = 3'b111; end
            18'b010101101011000100: begin rgb_reg = 3'b111; end
            18'b010101101011000101: begin rgb_reg = 3'b111; end
            18'b010101101011000110: begin rgb_reg = 3'b111; end
            18'b010101101011000111: begin rgb_reg = 3'b111; end
            18'b010101101011001100: begin rgb_reg = 3'b111; end
            18'b010101101011001101: begin rgb_reg = 3'b111; end
            18'b010101101011010000: begin rgb_reg = 3'b111; end
            18'b010101101011010001: begin rgb_reg = 3'b111; end
            18'b010101101011010010: begin rgb_reg = 3'b111; end
            18'b010101101011010011: begin rgb_reg = 3'b111; end
            18'b010101101011011010: begin rgb_reg = 3'b111; end
            18'b010101101011011011: begin rgb_reg = 3'b111; end
            18'b010101101011011100: begin rgb_reg = 3'b111; end
            18'b010101101011011101: begin rgb_reg = 3'b111; end
            18'b010101101011011110: begin rgb_reg = 3'b111; end
            18'b010101101011011111: begin rgb_reg = 3'b111; end
            18'b010101101011100100: begin rgb_reg = 3'b111; end
            18'b010101101011100101: begin rgb_reg = 3'b111; end
            18'b010101101011101000: begin rgb_reg = 3'b111; end
            18'b010101101011101001: begin rgb_reg = 3'b111; end
            18'b010101101011101010: begin rgb_reg = 3'b111; end
            18'b010101101011101011: begin rgb_reg = 3'b111; end
            18'b010101101011110000: begin rgb_reg = 3'b111; end
            18'b010101101011110001: begin rgb_reg = 3'b111; end
            18'b010101101011110100: begin rgb_reg = 3'b111; end
            18'b010101101011110101: begin rgb_reg = 3'b111; end
            18'b010101101011110110: begin rgb_reg = 3'b111; end
            18'b010101101011110111: begin rgb_reg = 3'b111; end
            18'b010101101011111110: begin rgb_reg = 3'b111; end
            18'b010101101011111111: begin rgb_reg = 3'b111; end
            18'b010101101100000000: begin rgb_reg = 3'b111; end
            18'b010101101100000001: begin rgb_reg = 3'b111; end
            18'b010101101100000010: begin rgb_reg = 3'b111; end
            18'b010101101100000011: begin rgb_reg = 3'b111; end
            18'b010101101100001010: begin rgb_reg = 3'b111; end
            18'b010101101100001011: begin rgb_reg = 3'b111; end
            18'b010101101100011110: begin rgb_reg = 3'b111; end
            18'b010101101100011111: begin rgb_reg = 3'b111; end
            18'b010101101100100000: begin rgb_reg = 3'b111; end
            18'b010101101100100001: begin rgb_reg = 3'b111; end
            18'b010101101100100010: begin rgb_reg = 3'b111; end
            18'b010101101100100011: begin rgb_reg = 3'b111; end
            18'b010101101100101010: begin rgb_reg = 3'b111; end
            18'b010101101100101011: begin rgb_reg = 3'b111; end
            18'b010101101100101100: begin rgb_reg = 3'b111; end
            18'b010101101100101101: begin rgb_reg = 3'b111; end
            18'b010101101100101110: begin rgb_reg = 3'b111; end
            18'b010101101100101111: begin rgb_reg = 3'b111; end
            18'b010101101100110110: begin rgb_reg = 3'b111; end
            18'b010101101100110111: begin rgb_reg = 3'b111; end
            18'b010101101100111000: begin rgb_reg = 3'b111; end
            18'b010101101100111001: begin rgb_reg = 3'b111; end
            18'b010101101100111010: begin rgb_reg = 3'b111; end
            18'b010101101100111011: begin rgb_reg = 3'b111; end
            18'b010101101101000000: begin rgb_reg = 3'b111; end
            18'b010101101101000001: begin rgb_reg = 3'b111; end
            18'b010101101101001000: begin rgb_reg = 3'b111; end
            18'b010101101101001001: begin rgb_reg = 3'b111; end
            18'b010101101101001010: begin rgb_reg = 3'b111; end
            18'b010101101101001011: begin rgb_reg = 3'b111; end
            18'b010101101101001100: begin rgb_reg = 3'b111; end
            18'b010101101101001101: begin rgb_reg = 3'b111; end
            18'b010101110010110100: begin rgb_reg = 3'b111; end
            18'b010101110010110101: begin rgb_reg = 3'b111; end
            18'b010101110010111100: begin rgb_reg = 3'b111; end
            18'b010101110010111101: begin rgb_reg = 3'b111; end
            18'b010101110011000000: begin rgb_reg = 3'b111; end
            18'b010101110011000001: begin rgb_reg = 3'b111; end
            18'b010101110011001000: begin rgb_reg = 3'b111; end
            18'b010101110011001001: begin rgb_reg = 3'b111; end
            18'b010101110011001100: begin rgb_reg = 3'b111; end
            18'b010101110011001101: begin rgb_reg = 3'b111; end
            18'b010101110011001110: begin rgb_reg = 3'b111; end
            18'b010101110011001111: begin rgb_reg = 3'b111; end
            18'b010101110011010100: begin rgb_reg = 3'b111; end
            18'b010101110011010101: begin rgb_reg = 3'b111; end
            18'b010101110011100000: begin rgb_reg = 3'b111; end
            18'b010101110011100001: begin rgb_reg = 3'b111; end
            18'b010101110011100100: begin rgb_reg = 3'b111; end
            18'b010101110011100101: begin rgb_reg = 3'b111; end
            18'b010101110011100110: begin rgb_reg = 3'b111; end
            18'b010101110011100111: begin rgb_reg = 3'b111; end
            18'b010101110011101100: begin rgb_reg = 3'b111; end
            18'b010101110011101101: begin rgb_reg = 3'b111; end
            18'b010101110011110000: begin rgb_reg = 3'b111; end
            18'b010101110011110001: begin rgb_reg = 3'b111; end
            18'b010101110011110010: begin rgb_reg = 3'b111; end
            18'b010101110011110011: begin rgb_reg = 3'b111; end
            18'b010101110011111000: begin rgb_reg = 3'b111; end
            18'b010101110011111001: begin rgb_reg = 3'b111; end
            18'b010101110100000100: begin rgb_reg = 3'b111; end
            18'b010101110100000101: begin rgb_reg = 3'b111; end
            18'b010101110100001010: begin rgb_reg = 3'b111; end
            18'b010101110100001011: begin rgb_reg = 3'b111; end
            18'b010101110100100100: begin rgb_reg = 3'b111; end
            18'b010101110100100101: begin rgb_reg = 3'b111; end
            18'b010101110100110000: begin rgb_reg = 3'b111; end
            18'b010101110100110001: begin rgb_reg = 3'b111; end
            18'b010101110100110100: begin rgb_reg = 3'b111; end
            18'b010101110100110101: begin rgb_reg = 3'b111; end
            18'b010101110100111100: begin rgb_reg = 3'b111; end
            18'b010101110100111101: begin rgb_reg = 3'b111; end
            18'b010101110101000000: begin rgb_reg = 3'b111; end
            18'b010101110101000001: begin rgb_reg = 3'b111; end
            18'b010101110101000110: begin rgb_reg = 3'b111; end
            18'b010101110101000111: begin rgb_reg = 3'b111; end
            18'b010101110101001110: begin rgb_reg = 3'b111; end
            18'b010101110101001111: begin rgb_reg = 3'b111; end
            18'b010101111010110100: begin rgb_reg = 3'b111; end
            18'b010101111010110101: begin rgb_reg = 3'b111; end
            18'b010101111010111100: begin rgb_reg = 3'b111; end
            18'b010101111010111101: begin rgb_reg = 3'b111; end
            18'b010101111011000000: begin rgb_reg = 3'b111; end
            18'b010101111011000001: begin rgb_reg = 3'b111; end
            18'b010101111011001000: begin rgb_reg = 3'b111; end
            18'b010101111011001001: begin rgb_reg = 3'b111; end
            18'b010101111011001100: begin rgb_reg = 3'b111; end
            18'b010101111011001101: begin rgb_reg = 3'b111; end
            18'b010101111011001110: begin rgb_reg = 3'b111; end
            18'b010101111011001111: begin rgb_reg = 3'b111; end
            18'b010101111011010100: begin rgb_reg = 3'b111; end
            18'b010101111011010101: begin rgb_reg = 3'b111; end
            18'b010101111011100000: begin rgb_reg = 3'b111; end
            18'b010101111011100001: begin rgb_reg = 3'b111; end
            18'b010101111011100100: begin rgb_reg = 3'b111; end
            18'b010101111011100101: begin rgb_reg = 3'b111; end
            18'b010101111011100110: begin rgb_reg = 3'b111; end
            18'b010101111011100111: begin rgb_reg = 3'b111; end
            18'b010101111011101100: begin rgb_reg = 3'b111; end
            18'b010101111011101101: begin rgb_reg = 3'b111; end
            18'b010101111011110000: begin rgb_reg = 3'b111; end
            18'b010101111011110001: begin rgb_reg = 3'b111; end
            18'b010101111011110010: begin rgb_reg = 3'b111; end
            18'b010101111011110011: begin rgb_reg = 3'b111; end
            18'b010101111011111000: begin rgb_reg = 3'b111; end
            18'b010101111011111001: begin rgb_reg = 3'b111; end
            18'b010101111100000100: begin rgb_reg = 3'b111; end
            18'b010101111100000101: begin rgb_reg = 3'b111; end
            18'b010101111100001010: begin rgb_reg = 3'b111; end
            18'b010101111100001011: begin rgb_reg = 3'b111; end
            18'b010101111100100100: begin rgb_reg = 3'b111; end
            18'b010101111100100101: begin rgb_reg = 3'b111; end
            18'b010101111100110000: begin rgb_reg = 3'b111; end
            18'b010101111100110001: begin rgb_reg = 3'b111; end
            18'b010101111100110100: begin rgb_reg = 3'b111; end
            18'b010101111100110101: begin rgb_reg = 3'b111; end
            18'b010101111100111100: begin rgb_reg = 3'b111; end
            18'b010101111100111101: begin rgb_reg = 3'b111; end
            18'b010101111101000000: begin rgb_reg = 3'b111; end
            18'b010101111101000001: begin rgb_reg = 3'b111; end
            18'b010101111101000110: begin rgb_reg = 3'b111; end
            18'b010101111101000111: begin rgb_reg = 3'b111; end
            18'b010101111101001110: begin rgb_reg = 3'b111; end
            18'b010101111101001111: begin rgb_reg = 3'b111; end
            18'b010110000010110100: begin rgb_reg = 3'b111; end
            18'b010110000010110101: begin rgb_reg = 3'b111; end
            18'b010110000010111000: begin rgb_reg = 3'b111; end
            18'b010110000010111001: begin rgb_reg = 3'b111; end
            18'b010110000010111100: begin rgb_reg = 3'b111; end
            18'b010110000010111101: begin rgb_reg = 3'b111; end
            18'b010110000011000000: begin rgb_reg = 3'b111; end
            18'b010110000011000001: begin rgb_reg = 3'b111; end
            18'b010110000011001000: begin rgb_reg = 3'b111; end
            18'b010110000011001001: begin rgb_reg = 3'b111; end
            18'b010110000011001100: begin rgb_reg = 3'b111; end
            18'b010110000011001101: begin rgb_reg = 3'b111; end
            18'b010110000011011010: begin rgb_reg = 3'b111; end
            18'b010110000011011011: begin rgb_reg = 3'b111; end
            18'b010110000011011100: begin rgb_reg = 3'b111; end
            18'b010110000011011101: begin rgb_reg = 3'b111; end
            18'b010110000011011110: begin rgb_reg = 3'b111; end
            18'b010110000011011111: begin rgb_reg = 3'b111; end
            18'b010110000011100000: begin rgb_reg = 3'b111; end
            18'b010110000011100001: begin rgb_reg = 3'b111; end
            18'b010110000011100100: begin rgb_reg = 3'b111; end
            18'b010110000011100101: begin rgb_reg = 3'b111; end
            18'b010110000011101100: begin rgb_reg = 3'b111; end
            18'b010110000011101101: begin rgb_reg = 3'b111; end
            18'b010110000011110000: begin rgb_reg = 3'b111; end
            18'b010110000011110001: begin rgb_reg = 3'b111; end
            18'b010110000011111110: begin rgb_reg = 3'b111; end
            18'b010110000011111111: begin rgb_reg = 3'b111; end
            18'b010110000100000000: begin rgb_reg = 3'b111; end
            18'b010110000100000001: begin rgb_reg = 3'b111; end
            18'b010110000100000010: begin rgb_reg = 3'b111; end
            18'b010110000100000011: begin rgb_reg = 3'b111; end
            18'b010110000100000100: begin rgb_reg = 3'b111; end
            18'b010110000100000101: begin rgb_reg = 3'b111; end
            18'b010110000100001010: begin rgb_reg = 3'b111; end
            18'b010110000100001011: begin rgb_reg = 3'b111; end
            18'b010110000100100100: begin rgb_reg = 3'b111; end
            18'b010110000100100101: begin rgb_reg = 3'b111; end
            18'b010110000100101010: begin rgb_reg = 3'b111; end
            18'b010110000100101011: begin rgb_reg = 3'b111; end
            18'b010110000100101100: begin rgb_reg = 3'b111; end
            18'b010110000100101101: begin rgb_reg = 3'b111; end
            18'b010110000100101110: begin rgb_reg = 3'b111; end
            18'b010110000100101111: begin rgb_reg = 3'b111; end
            18'b010110000100110000: begin rgb_reg = 3'b111; end
            18'b010110000100110001: begin rgb_reg = 3'b111; end
            18'b010110000100110100: begin rgb_reg = 3'b111; end
            18'b010110000100110101: begin rgb_reg = 3'b111; end
            18'b010110000100110110: begin rgb_reg = 3'b111; end
            18'b010110000100110111: begin rgb_reg = 3'b111; end
            18'b010110000100111000: begin rgb_reg = 3'b111; end
            18'b010110000100111001: begin rgb_reg = 3'b111; end
            18'b010110000100111010: begin rgb_reg = 3'b111; end
            18'b010110000100111011: begin rgb_reg = 3'b111; end
            18'b010110000100111100: begin rgb_reg = 3'b111; end
            18'b010110000100111101: begin rgb_reg = 3'b111; end
            18'b010110000101000000: begin rgb_reg = 3'b111; end
            18'b010110000101000001: begin rgb_reg = 3'b111; end
            18'b010110000101000110: begin rgb_reg = 3'b111; end
            18'b010110000101000111: begin rgb_reg = 3'b111; end
            18'b010110000101001110: begin rgb_reg = 3'b111; end
            18'b010110000101001111: begin rgb_reg = 3'b111; end
            18'b010110001010110100: begin rgb_reg = 3'b111; end
            18'b010110001010110101: begin rgb_reg = 3'b111; end
            18'b010110001010111000: begin rgb_reg = 3'b111; end
            18'b010110001010111001: begin rgb_reg = 3'b111; end
            18'b010110001010111100: begin rgb_reg = 3'b111; end
            18'b010110001010111101: begin rgb_reg = 3'b111; end
            18'b010110001011000000: begin rgb_reg = 3'b111; end
            18'b010110001011000001: begin rgb_reg = 3'b111; end
            18'b010110001011001000: begin rgb_reg = 3'b111; end
            18'b010110001011001001: begin rgb_reg = 3'b111; end
            18'b010110001011001100: begin rgb_reg = 3'b111; end
            18'b010110001011001101: begin rgb_reg = 3'b111; end
            18'b010110001011011010: begin rgb_reg = 3'b111; end
            18'b010110001011011011: begin rgb_reg = 3'b111; end
            18'b010110001011011100: begin rgb_reg = 3'b111; end
            18'b010110001011011101: begin rgb_reg = 3'b111; end
            18'b010110001011011110: begin rgb_reg = 3'b111; end
            18'b010110001011011111: begin rgb_reg = 3'b111; end
            18'b010110001011100000: begin rgb_reg = 3'b111; end
            18'b010110001011100001: begin rgb_reg = 3'b111; end
            18'b010110001011100100: begin rgb_reg = 3'b111; end
            18'b010110001011100101: begin rgb_reg = 3'b111; end
            18'b010110001011101100: begin rgb_reg = 3'b111; end
            18'b010110001011101101: begin rgb_reg = 3'b111; end
            18'b010110001011110000: begin rgb_reg = 3'b111; end
            18'b010110001011110001: begin rgb_reg = 3'b111; end
            18'b010110001011111110: begin rgb_reg = 3'b111; end
            18'b010110001011111111: begin rgb_reg = 3'b111; end
            18'b010110001100000000: begin rgb_reg = 3'b111; end
            18'b010110001100000001: begin rgb_reg = 3'b111; end
            18'b010110001100000010: begin rgb_reg = 3'b111; end
            18'b010110001100000011: begin rgb_reg = 3'b111; end
            18'b010110001100000100: begin rgb_reg = 3'b111; end
            18'b010110001100000101: begin rgb_reg = 3'b111; end
            18'b010110001100001010: begin rgb_reg = 3'b111; end
            18'b010110001100001011: begin rgb_reg = 3'b111; end
            18'b010110001100100100: begin rgb_reg = 3'b111; end
            18'b010110001100100101: begin rgb_reg = 3'b111; end
            18'b010110001100101010: begin rgb_reg = 3'b111; end
            18'b010110001100101011: begin rgb_reg = 3'b111; end
            18'b010110001100101100: begin rgb_reg = 3'b111; end
            18'b010110001100101101: begin rgb_reg = 3'b111; end
            18'b010110001100101110: begin rgb_reg = 3'b111; end
            18'b010110001100101111: begin rgb_reg = 3'b111; end
            18'b010110001100110000: begin rgb_reg = 3'b111; end
            18'b010110001100110001: begin rgb_reg = 3'b111; end
            18'b010110001100110100: begin rgb_reg = 3'b111; end
            18'b010110001100110101: begin rgb_reg = 3'b111; end
            18'b010110001100110110: begin rgb_reg = 3'b111; end
            18'b010110001100110111: begin rgb_reg = 3'b111; end
            18'b010110001100111000: begin rgb_reg = 3'b111; end
            18'b010110001100111001: begin rgb_reg = 3'b111; end
            18'b010110001100111010: begin rgb_reg = 3'b111; end
            18'b010110001100111011: begin rgb_reg = 3'b111; end
            18'b010110001100111100: begin rgb_reg = 3'b111; end
            18'b010110001100111101: begin rgb_reg = 3'b111; end
            18'b010110001101000000: begin rgb_reg = 3'b111; end
            18'b010110001101000001: begin rgb_reg = 3'b111; end
            18'b010110001101000110: begin rgb_reg = 3'b111; end
            18'b010110001101000111: begin rgb_reg = 3'b111; end
            18'b010110001101001110: begin rgb_reg = 3'b111; end
            18'b010110001101001111: begin rgb_reg = 3'b111; end
            18'b010110010010110100: begin rgb_reg = 3'b111; end
            18'b010110010010110101: begin rgb_reg = 3'b111; end
            18'b010110010010110110: begin rgb_reg = 3'b111; end
            18'b010110010010110111: begin rgb_reg = 3'b111; end
            18'b010110010010111010: begin rgb_reg = 3'b111; end
            18'b010110010010111011: begin rgb_reg = 3'b111; end
            18'b010110010010111100: begin rgb_reg = 3'b111; end
            18'b010110010010111101: begin rgb_reg = 3'b111; end
            18'b010110010011000000: begin rgb_reg = 3'b111; end
            18'b010110010011000001: begin rgb_reg = 3'b111; end
            18'b010110010011001000: begin rgb_reg = 3'b111; end
            18'b010110010011001001: begin rgb_reg = 3'b111; end
            18'b010110010011001100: begin rgb_reg = 3'b111; end
            18'b010110010011001101: begin rgb_reg = 3'b111; end
            18'b010110010011011000: begin rgb_reg = 3'b111; end
            18'b010110010011011001: begin rgb_reg = 3'b111; end
            18'b010110010011100000: begin rgb_reg = 3'b111; end
            18'b010110010011100001: begin rgb_reg = 3'b111; end
            18'b010110010011100100: begin rgb_reg = 3'b111; end
            18'b010110010011100101: begin rgb_reg = 3'b111; end
            18'b010110010011100110: begin rgb_reg = 3'b111; end
            18'b010110010011100111: begin rgb_reg = 3'b111; end
            18'b010110010011101000: begin rgb_reg = 3'b111; end
            18'b010110010011101001: begin rgb_reg = 3'b111; end
            18'b010110010011101010: begin rgb_reg = 3'b111; end
            18'b010110010011101011: begin rgb_reg = 3'b111; end
            18'b010110010011110000: begin rgb_reg = 3'b111; end
            18'b010110010011110001: begin rgb_reg = 3'b111; end
            18'b010110010011111100: begin rgb_reg = 3'b111; end
            18'b010110010011111101: begin rgb_reg = 3'b111; end
            18'b010110010100000100: begin rgb_reg = 3'b111; end
            18'b010110010100000101: begin rgb_reg = 3'b111; end
            18'b010110010100001010: begin rgb_reg = 3'b111; end
            18'b010110010100001011: begin rgb_reg = 3'b111; end
            18'b010110010100011100: begin rgb_reg = 3'b111; end
            18'b010110010100011101: begin rgb_reg = 3'b111; end
            18'b010110010100100100: begin rgb_reg = 3'b111; end
            18'b010110010100100101: begin rgb_reg = 3'b111; end
            18'b010110010100101000: begin rgb_reg = 3'b111; end
            18'b010110010100101001: begin rgb_reg = 3'b111; end
            18'b010110010100110000: begin rgb_reg = 3'b111; end
            18'b010110010100110001: begin rgb_reg = 3'b111; end
            18'b010110010100110100: begin rgb_reg = 3'b111; end
            18'b010110010100110101: begin rgb_reg = 3'b111; end
            18'b010110010101000000: begin rgb_reg = 3'b111; end
            18'b010110010101000001: begin rgb_reg = 3'b111; end
            18'b010110010101000110: begin rgb_reg = 3'b111; end
            18'b010110010101000111: begin rgb_reg = 3'b111; end
            18'b010110010101001110: begin rgb_reg = 3'b111; end
            18'b010110010101001111: begin rgb_reg = 3'b111; end
            18'b010110011010110100: begin rgb_reg = 3'b111; end
            18'b010110011010110101: begin rgb_reg = 3'b111; end
            18'b010110011010110110: begin rgb_reg = 3'b111; end
            18'b010110011010110111: begin rgb_reg = 3'b111; end
            18'b010110011010111010: begin rgb_reg = 3'b111; end
            18'b010110011010111011: begin rgb_reg = 3'b111; end
            18'b010110011010111100: begin rgb_reg = 3'b111; end
            18'b010110011010111101: begin rgb_reg = 3'b111; end
            18'b010110011011000000: begin rgb_reg = 3'b111; end
            18'b010110011011000001: begin rgb_reg = 3'b111; end
            18'b010110011011001000: begin rgb_reg = 3'b111; end
            18'b010110011011001001: begin rgb_reg = 3'b111; end
            18'b010110011011001100: begin rgb_reg = 3'b111; end
            18'b010110011011001101: begin rgb_reg = 3'b111; end
            18'b010110011011011000: begin rgb_reg = 3'b111; end
            18'b010110011011011001: begin rgb_reg = 3'b111; end
            18'b010110011011100000: begin rgb_reg = 3'b111; end
            18'b010110011011100001: begin rgb_reg = 3'b111; end
            18'b010110011011100100: begin rgb_reg = 3'b111; end
            18'b010110011011100101: begin rgb_reg = 3'b111; end
            18'b010110011011100110: begin rgb_reg = 3'b111; end
            18'b010110011011100111: begin rgb_reg = 3'b111; end
            18'b010110011011101000: begin rgb_reg = 3'b111; end
            18'b010110011011101001: begin rgb_reg = 3'b111; end
            18'b010110011011101010: begin rgb_reg = 3'b111; end
            18'b010110011011101011: begin rgb_reg = 3'b111; end
            18'b010110011011110000: begin rgb_reg = 3'b111; end
            18'b010110011011110001: begin rgb_reg = 3'b111; end
            18'b010110011011111100: begin rgb_reg = 3'b111; end
            18'b010110011011111101: begin rgb_reg = 3'b111; end
            18'b010110011100000100: begin rgb_reg = 3'b111; end
            18'b010110011100000101: begin rgb_reg = 3'b111; end
            18'b010110011100001010: begin rgb_reg = 3'b111; end
            18'b010110011100001011: begin rgb_reg = 3'b111; end
            18'b010110011100011100: begin rgb_reg = 3'b111; end
            18'b010110011100011101: begin rgb_reg = 3'b111; end
            18'b010110011100100100: begin rgb_reg = 3'b111; end
            18'b010110011100100101: begin rgb_reg = 3'b111; end
            18'b010110011100101000: begin rgb_reg = 3'b111; end
            18'b010110011100101001: begin rgb_reg = 3'b111; end
            18'b010110011100110000: begin rgb_reg = 3'b111; end
            18'b010110011100110001: begin rgb_reg = 3'b111; end
            18'b010110011100110100: begin rgb_reg = 3'b111; end
            18'b010110011100110101: begin rgb_reg = 3'b111; end
            18'b010110011101000000: begin rgb_reg = 3'b111; end
            18'b010110011101000001: begin rgb_reg = 3'b111; end
            18'b010110011101000110: begin rgb_reg = 3'b111; end
            18'b010110011101000111: begin rgb_reg = 3'b111; end
            18'b010110011101001110: begin rgb_reg = 3'b111; end
            18'b010110011101001111: begin rgb_reg = 3'b111; end
            18'b010110100010110100: begin rgb_reg = 3'b111; end
            18'b010110100010110101: begin rgb_reg = 3'b111; end
            18'b010110100010111100: begin rgb_reg = 3'b111; end
            18'b010110100010111101: begin rgb_reg = 3'b111; end
            18'b010110100011000010: begin rgb_reg = 3'b111; end
            18'b010110100011000011: begin rgb_reg = 3'b111; end
            18'b010110100011000100: begin rgb_reg = 3'b111; end
            18'b010110100011000101: begin rgb_reg = 3'b111; end
            18'b010110100011000110: begin rgb_reg = 3'b111; end
            18'b010110100011000111: begin rgb_reg = 3'b111; end
            18'b010110100011001100: begin rgb_reg = 3'b111; end
            18'b010110100011001101: begin rgb_reg = 3'b111; end
            18'b010110100011011010: begin rgb_reg = 3'b111; end
            18'b010110100011011011: begin rgb_reg = 3'b111; end
            18'b010110100011011100: begin rgb_reg = 3'b111; end
            18'b010110100011011101: begin rgb_reg = 3'b111; end
            18'b010110100011011110: begin rgb_reg = 3'b111; end
            18'b010110100011011111: begin rgb_reg = 3'b111; end
            18'b010110100011100000: begin rgb_reg = 3'b111; end
            18'b010110100011100001: begin rgb_reg = 3'b111; end
            18'b010110100011100100: begin rgb_reg = 3'b111; end
            18'b010110100011100101: begin rgb_reg = 3'b111; end
            18'b010110100011110000: begin rgb_reg = 3'b111; end
            18'b010110100011110001: begin rgb_reg = 3'b111; end
            18'b010110100011111110: begin rgb_reg = 3'b111; end
            18'b010110100011111111: begin rgb_reg = 3'b111; end
            18'b010110100100000000: begin rgb_reg = 3'b111; end
            18'b010110100100000001: begin rgb_reg = 3'b111; end
            18'b010110100100000010: begin rgb_reg = 3'b111; end
            18'b010110100100000011: begin rgb_reg = 3'b111; end
            18'b010110100100000100: begin rgb_reg = 3'b111; end
            18'b010110100100000101: begin rgb_reg = 3'b111; end
            18'b010110100100001100: begin rgb_reg = 3'b111; end
            18'b010110100100001101: begin rgb_reg = 3'b111; end
            18'b010110100100011110: begin rgb_reg = 3'b111; end
            18'b010110100100011111: begin rgb_reg = 3'b111; end
            18'b010110100100100000: begin rgb_reg = 3'b111; end
            18'b010110100100100001: begin rgb_reg = 3'b111; end
            18'b010110100100100010: begin rgb_reg = 3'b111; end
            18'b010110100100100011: begin rgb_reg = 3'b111; end
            18'b010110100100101010: begin rgb_reg = 3'b111; end
            18'b010110100100101011: begin rgb_reg = 3'b111; end
            18'b010110100100101100: begin rgb_reg = 3'b111; end
            18'b010110100100101101: begin rgb_reg = 3'b111; end
            18'b010110100100101110: begin rgb_reg = 3'b111; end
            18'b010110100100101111: begin rgb_reg = 3'b111; end
            18'b010110100100110000: begin rgb_reg = 3'b111; end
            18'b010110100100110001: begin rgb_reg = 3'b111; end
            18'b010110100100110110: begin rgb_reg = 3'b111; end
            18'b010110100100110111: begin rgb_reg = 3'b111; end
            18'b010110100100111000: begin rgb_reg = 3'b111; end
            18'b010110100100111001: begin rgb_reg = 3'b111; end
            18'b010110100100111010: begin rgb_reg = 3'b111; end
            18'b010110100100111011: begin rgb_reg = 3'b111; end
            18'b010110100100111100: begin rgb_reg = 3'b111; end
            18'b010110100100111101: begin rgb_reg = 3'b111; end
            18'b010110100101000010: begin rgb_reg = 3'b111; end
            18'b010110100101000011: begin rgb_reg = 3'b111; end
            18'b010110100101001000: begin rgb_reg = 3'b111; end
            18'b010110100101001001: begin rgb_reg = 3'b111; end
            18'b010110100101001010: begin rgb_reg = 3'b111; end
            18'b010110100101001011: begin rgb_reg = 3'b111; end
            18'b010110100101001100: begin rgb_reg = 3'b111; end
            18'b010110100101001101: begin rgb_reg = 3'b111; end
            18'b010110101010110100: begin rgb_reg = 3'b111; end
            18'b010110101010110101: begin rgb_reg = 3'b111; end
            18'b010110101010111100: begin rgb_reg = 3'b111; end
            18'b010110101010111101: begin rgb_reg = 3'b111; end
            18'b010110101011000010: begin rgb_reg = 3'b111; end
            18'b010110101011000011: begin rgb_reg = 3'b111; end
            18'b010110101011000100: begin rgb_reg = 3'b111; end
            18'b010110101011000101: begin rgb_reg = 3'b111; end
            18'b010110101011000110: begin rgb_reg = 3'b111; end
            18'b010110101011000111: begin rgb_reg = 3'b111; end
            18'b010110101011001100: begin rgb_reg = 3'b111; end
            18'b010110101011001101: begin rgb_reg = 3'b111; end
            18'b010110101011011010: begin rgb_reg = 3'b111; end
            18'b010110101011011011: begin rgb_reg = 3'b111; end
            18'b010110101011011100: begin rgb_reg = 3'b111; end
            18'b010110101011011101: begin rgb_reg = 3'b111; end
            18'b010110101011011110: begin rgb_reg = 3'b111; end
            18'b010110101011011111: begin rgb_reg = 3'b111; end
            18'b010110101011100000: begin rgb_reg = 3'b111; end
            18'b010110101011100001: begin rgb_reg = 3'b111; end
            18'b010110101011100100: begin rgb_reg = 3'b111; end
            18'b010110101011100101: begin rgb_reg = 3'b111; end
            18'b010110101011110000: begin rgb_reg = 3'b111; end
            18'b010110101011110001: begin rgb_reg = 3'b111; end
            18'b010110101011111110: begin rgb_reg = 3'b111; end
            18'b010110101011111111: begin rgb_reg = 3'b111; end
            18'b010110101100000000: begin rgb_reg = 3'b111; end
            18'b010110101100000001: begin rgb_reg = 3'b111; end
            18'b010110101100000010: begin rgb_reg = 3'b111; end
            18'b010110101100000011: begin rgb_reg = 3'b111; end
            18'b010110101100000100: begin rgb_reg = 3'b111; end
            18'b010110101100000101: begin rgb_reg = 3'b111; end
            18'b010110101100001100: begin rgb_reg = 3'b111; end
            18'b010110101100001101: begin rgb_reg = 3'b111; end
            18'b010110101100011110: begin rgb_reg = 3'b111; end
            18'b010110101100011111: begin rgb_reg = 3'b111; end
            18'b010110101100100000: begin rgb_reg = 3'b111; end
            18'b010110101100100001: begin rgb_reg = 3'b111; end
            18'b010110101100100010: begin rgb_reg = 3'b111; end
            18'b010110101100100011: begin rgb_reg = 3'b111; end
            18'b010110101100101010: begin rgb_reg = 3'b111; end
            18'b010110101100101011: begin rgb_reg = 3'b111; end
            18'b010110101100101100: begin rgb_reg = 3'b111; end
            18'b010110101100101101: begin rgb_reg = 3'b111; end
            18'b010110101100101110: begin rgb_reg = 3'b111; end
            18'b010110101100101111: begin rgb_reg = 3'b111; end
            18'b010110101100110000: begin rgb_reg = 3'b111; end
            18'b010110101100110001: begin rgb_reg = 3'b111; end
            18'b010110101100110110: begin rgb_reg = 3'b111; end
            18'b010110101100110111: begin rgb_reg = 3'b111; end
            18'b010110101100111000: begin rgb_reg = 3'b111; end
            18'b010110101100111001: begin rgb_reg = 3'b111; end
            18'b010110101100111010: begin rgb_reg = 3'b111; end
            18'b010110101100111011: begin rgb_reg = 3'b111; end
            18'b010110101100111100: begin rgb_reg = 3'b111; end
            18'b010110101100111101: begin rgb_reg = 3'b111; end
            18'b010110101101000010: begin rgb_reg = 3'b111; end
            18'b010110101101000011: begin rgb_reg = 3'b111; end
            18'b010110101101001000: begin rgb_reg = 3'b111; end
            18'b010110101101001001: begin rgb_reg = 3'b111; end
            18'b010110101101001010: begin rgb_reg = 3'b111; end
            18'b010110101101001011: begin rgb_reg = 3'b111; end
            18'b010110101101001100: begin rgb_reg = 3'b111; end
            18'b010110101101001101: begin rgb_reg = 3'b111; end
            18'b010110110011100100: begin rgb_reg = 3'b111; end
            18'b010110110011100101: begin rgb_reg = 3'b111; end
            18'b010110111011100100: begin rgb_reg = 3'b111; end
            18'b010110111011100101: begin rgb_reg = 3'b111; end
            18'b011001011011000010: begin rgb_reg = 3'b111; end
            18'b011001011011000011: begin rgb_reg = 3'b111; end
            18'b011001011011000100: begin rgb_reg = 3'b111; end
            18'b011001011011000101: begin rgb_reg = 3'b111; end
            18'b011001011011000110: begin rgb_reg = 3'b111; end
            18'b011001011011001101: begin rgb_reg = 3'b111; end
            18'b011001011011001110: begin rgb_reg = 3'b111; end
            18'b011001011011001111: begin rgb_reg = 3'b111; end
            18'b011001011011010000: begin rgb_reg = 3'b111; end
            18'b011001011011010001: begin rgb_reg = 3'b111; end
            18'b011001011011010010: begin rgb_reg = 3'b111; end
            18'b011001011011010011: begin rgb_reg = 3'b111; end
            18'b011001011011011011: begin rgb_reg = 3'b111; end
            18'b011001011011011100: begin rgb_reg = 3'b111; end
            18'b011001011011011101: begin rgb_reg = 3'b111; end
            18'b011001011011011110: begin rgb_reg = 3'b111; end
            18'b011001011011011111: begin rgb_reg = 3'b111; end
            18'b011001011011100000: begin rgb_reg = 3'b111; end
            18'b011001011011100001: begin rgb_reg = 3'b111; end
            18'b011001011011101011: begin rgb_reg = 3'b111; end
            18'b011001011011101100: begin rgb_reg = 3'b111; end
            18'b011001011011110110: begin rgb_reg = 3'b111; end
            18'b011001011011110111: begin rgb_reg = 3'b111; end
            18'b011001011011111000: begin rgb_reg = 3'b111; end
            18'b011001011011111001: begin rgb_reg = 3'b111; end
            18'b011001011011111010: begin rgb_reg = 3'b111; end
            18'b011001011011111011: begin rgb_reg = 3'b111; end
            18'b011001011011111100: begin rgb_reg = 3'b111; end
            18'b011001011100000110: begin rgb_reg = 3'b111; end
            18'b011001011100000111: begin rgb_reg = 3'b111; end
            18'b011001011100001000: begin rgb_reg = 3'b111; end
            18'b011001011100001001: begin rgb_reg = 3'b111; end
            18'b011001011100010011: begin rgb_reg = 3'b111; end
            18'b011001011100010100: begin rgb_reg = 3'b111; end
            18'b011001011100010101: begin rgb_reg = 3'b111; end
            18'b011001011100011110: begin rgb_reg = 3'b111; end
            18'b011001011100011111: begin rgb_reg = 3'b111; end
            18'b011001011100100000: begin rgb_reg = 3'b111; end
            18'b011001011100100001: begin rgb_reg = 3'b111; end
            18'b011001011100100010: begin rgb_reg = 3'b111; end
            18'b011001011100100011: begin rgb_reg = 3'b111; end
            18'b011001011100100100: begin rgb_reg = 3'b111; end
            18'b011001011100101100: begin rgb_reg = 3'b111; end
            18'b011001011100101101: begin rgb_reg = 3'b111; end
            18'b011001011100101110: begin rgb_reg = 3'b111; end
            18'b011001011100101111: begin rgb_reg = 3'b111; end
            18'b011001011100110000: begin rgb_reg = 3'b111; end
            18'b011001011100110001: begin rgb_reg = 3'b111; end
            18'b011001011100110010: begin rgb_reg = 3'b111; end
            18'b011001011100111100: begin rgb_reg = 3'b111; end
            18'b011001011100111101: begin rgb_reg = 3'b111; end
            18'b011001100011000010: begin rgb_reg = 3'b111; end
            18'b011001100011000011: begin rgb_reg = 3'b111; end
            18'b011001100011000100: begin rgb_reg = 3'b111; end
            18'b011001100011000101: begin rgb_reg = 3'b111; end
            18'b011001100011000110: begin rgb_reg = 3'b111; end
            18'b011001100011001101: begin rgb_reg = 3'b111; end
            18'b011001100011001110: begin rgb_reg = 3'b111; end
            18'b011001100011001111: begin rgb_reg = 3'b111; end
            18'b011001100011010000: begin rgb_reg = 3'b111; end
            18'b011001100011010001: begin rgb_reg = 3'b111; end
            18'b011001100011010010: begin rgb_reg = 3'b111; end
            18'b011001100011010011: begin rgb_reg = 3'b111; end
            18'b011001100011011011: begin rgb_reg = 3'b111; end
            18'b011001100011011100: begin rgb_reg = 3'b111; end
            18'b011001100011011101: begin rgb_reg = 3'b111; end
            18'b011001100011011110: begin rgb_reg = 3'b111; end
            18'b011001100011011111: begin rgb_reg = 3'b111; end
            18'b011001100011100000: begin rgb_reg = 3'b111; end
            18'b011001100011100001: begin rgb_reg = 3'b111; end
            18'b011001100011101011: begin rgb_reg = 3'b111; end
            18'b011001100011101100: begin rgb_reg = 3'b111; end
            18'b011001100011110110: begin rgb_reg = 3'b111; end
            18'b011001100011110111: begin rgb_reg = 3'b111; end
            18'b011001100011111000: begin rgb_reg = 3'b111; end
            18'b011001100011111001: begin rgb_reg = 3'b111; end
            18'b011001100011111010: begin rgb_reg = 3'b111; end
            18'b011001100011111011: begin rgb_reg = 3'b111; end
            18'b011001100011111100: begin rgb_reg = 3'b111; end
            18'b011001100100000110: begin rgb_reg = 3'b111; end
            18'b011001100100000111: begin rgb_reg = 3'b111; end
            18'b011001100100001000: begin rgb_reg = 3'b111; end
            18'b011001100100001001: begin rgb_reg = 3'b111; end
            18'b011001100100010011: begin rgb_reg = 3'b111; end
            18'b011001100100010100: begin rgb_reg = 3'b111; end
            18'b011001100100010101: begin rgb_reg = 3'b111; end
            18'b011001100100011110: begin rgb_reg = 3'b111; end
            18'b011001100100011111: begin rgb_reg = 3'b111; end
            18'b011001100100100000: begin rgb_reg = 3'b111; end
            18'b011001100100100001: begin rgb_reg = 3'b111; end
            18'b011001100100100010: begin rgb_reg = 3'b111; end
            18'b011001100100100011: begin rgb_reg = 3'b111; end
            18'b011001100100100100: begin rgb_reg = 3'b111; end
            18'b011001100100101100: begin rgb_reg = 3'b111; end
            18'b011001100100101101: begin rgb_reg = 3'b111; end
            18'b011001100100101110: begin rgb_reg = 3'b111; end
            18'b011001100100101111: begin rgb_reg = 3'b111; end
            18'b011001100100110000: begin rgb_reg = 3'b111; end
            18'b011001100100110001: begin rgb_reg = 3'b111; end
            18'b011001100100110010: begin rgb_reg = 3'b111; end
            18'b011001100100111100: begin rgb_reg = 3'b111; end
            18'b011001100100111101: begin rgb_reg = 3'b111; end
            18'b011001101011000000: begin rgb_reg = 3'b111; end
            18'b011001101011000001: begin rgb_reg = 3'b111; end
            18'b011001101011001011: begin rgb_reg = 3'b111; end
            18'b011001101011001100: begin rgb_reg = 3'b111; end
            18'b011001101011001101: begin rgb_reg = 3'b111; end
            18'b011001101011010100: begin rgb_reg = 3'b111; end
            18'b011001101011010101: begin rgb_reg = 3'b111; end
            18'b011001101011011001: begin rgb_reg = 3'b111; end
            18'b011001101011011010: begin rgb_reg = 3'b111; end
            18'b011001101011100010: begin rgb_reg = 3'b111; end
            18'b011001101011100011: begin rgb_reg = 3'b111; end
            18'b011001101011101001: begin rgb_reg = 3'b111; end
            18'b011001101011101010: begin rgb_reg = 3'b111; end
            18'b011001101011101011: begin rgb_reg = 3'b111; end
            18'b011001101011101100: begin rgb_reg = 3'b111; end
            18'b011001101011110100: begin rgb_reg = 3'b111; end
            18'b011001101011110101: begin rgb_reg = 3'b111; end
            18'b011001101011111101: begin rgb_reg = 3'b111; end
            18'b011001101011111110: begin rgb_reg = 3'b111; end
            18'b011001101100000100: begin rgb_reg = 3'b111; end
            18'b011001101100000101: begin rgb_reg = 3'b111; end
            18'b011001101100010001: begin rgb_reg = 3'b111; end
            18'b011001101100010010: begin rgb_reg = 3'b111; end
            18'b011001101100010011: begin rgb_reg = 3'b111; end
            18'b011001101100010100: begin rgb_reg = 3'b111; end
            18'b011001101100010101: begin rgb_reg = 3'b111; end
            18'b011001101100011100: begin rgb_reg = 3'b111; end
            18'b011001101100011101: begin rgb_reg = 3'b111; end
            18'b011001101100011110: begin rgb_reg = 3'b111; end
            18'b011001101100100101: begin rgb_reg = 3'b111; end
            18'b011001101100100110: begin rgb_reg = 3'b111; end
            18'b011001101100101010: begin rgb_reg = 3'b111; end
            18'b011001101100101011: begin rgb_reg = 3'b111; end
            18'b011001101100110011: begin rgb_reg = 3'b111; end
            18'b011001101100110100: begin rgb_reg = 3'b111; end
            18'b011001101100111010: begin rgb_reg = 3'b111; end
            18'b011001101100111011: begin rgb_reg = 3'b111; end
            18'b011001101100111100: begin rgb_reg = 3'b111; end
            18'b011001101100111101: begin rgb_reg = 3'b111; end
            18'b011001110011000000: begin rgb_reg = 3'b111; end
            18'b011001110011000001: begin rgb_reg = 3'b111; end
            18'b011001110011001011: begin rgb_reg = 3'b111; end
            18'b011001110011001100: begin rgb_reg = 3'b111; end
            18'b011001110011001101: begin rgb_reg = 3'b111; end
            18'b011001110011010100: begin rgb_reg = 3'b111; end
            18'b011001110011010101: begin rgb_reg = 3'b111; end
            18'b011001110011010110: begin rgb_reg = 3'b111; end
            18'b011001110011011001: begin rgb_reg = 3'b111; end
            18'b011001110011011010: begin rgb_reg = 3'b111; end
            18'b011001110011100010: begin rgb_reg = 3'b111; end
            18'b011001110011100011: begin rgb_reg = 3'b111; end
            18'b011001110011101000: begin rgb_reg = 3'b111; end
            18'b011001110011101001: begin rgb_reg = 3'b111; end
            18'b011001110011101010: begin rgb_reg = 3'b111; end
            18'b011001110011101011: begin rgb_reg = 3'b111; end
            18'b011001110011101100: begin rgb_reg = 3'b111; end
            18'b011001110011110100: begin rgb_reg = 3'b111; end
            18'b011001110011110101: begin rgb_reg = 3'b111; end
            18'b011001110011111101: begin rgb_reg = 3'b111; end
            18'b011001110011111110: begin rgb_reg = 3'b111; end
            18'b011001110100000011: begin rgb_reg = 3'b111; end
            18'b011001110100000100: begin rgb_reg = 3'b111; end
            18'b011001110100000101: begin rgb_reg = 3'b111; end
            18'b011001110100010001: begin rgb_reg = 3'b111; end
            18'b011001110100010010: begin rgb_reg = 3'b111; end
            18'b011001110100010011: begin rgb_reg = 3'b111; end
            18'b011001110100010100: begin rgb_reg = 3'b111; end
            18'b011001110100010101: begin rgb_reg = 3'b111; end
            18'b011001110100011100: begin rgb_reg = 3'b111; end
            18'b011001110100011101: begin rgb_reg = 3'b111; end
            18'b011001110100011110: begin rgb_reg = 3'b111; end
            18'b011001110100100101: begin rgb_reg = 3'b111; end
            18'b011001110100100110: begin rgb_reg = 3'b111; end
            18'b011001110100100111: begin rgb_reg = 3'b111; end
            18'b011001110100101010: begin rgb_reg = 3'b111; end
            18'b011001110100101011: begin rgb_reg = 3'b111; end
            18'b011001110100110011: begin rgb_reg = 3'b111; end
            18'b011001110100110100: begin rgb_reg = 3'b111; end
            18'b011001110100111001: begin rgb_reg = 3'b111; end
            18'b011001110100111010: begin rgb_reg = 3'b111; end
            18'b011001110100111011: begin rgb_reg = 3'b111; end
            18'b011001110100111100: begin rgb_reg = 3'b111; end
            18'b011001110100111101: begin rgb_reg = 3'b111; end
            18'b011001111010111110: begin rgb_reg = 3'b111; end
            18'b011001111010111111: begin rgb_reg = 3'b111; end
            18'b011001111011000000: begin rgb_reg = 3'b111; end
            18'b011001111011000001: begin rgb_reg = 3'b111; end
            18'b011001111011001011: begin rgb_reg = 3'b111; end
            18'b011001111011001100: begin rgb_reg = 3'b111; end
            18'b011001111011001101: begin rgb_reg = 3'b111; end
            18'b011001111011010010: begin rgb_reg = 3'b111; end
            18'b011001111011010011: begin rgb_reg = 3'b111; end
            18'b011001111011010100: begin rgb_reg = 3'b111; end
            18'b011001111011010101: begin rgb_reg = 3'b111; end
            18'b011001111011010110: begin rgb_reg = 3'b111; end
            18'b011001111011011001: begin rgb_reg = 3'b111; end
            18'b011001111011011010: begin rgb_reg = 3'b111; end
            18'b011001111011100010: begin rgb_reg = 3'b111; end
            18'b011001111011100011: begin rgb_reg = 3'b111; end
            18'b011001111011101001: begin rgb_reg = 3'b111; end
            18'b011001111011101010: begin rgb_reg = 3'b111; end
            18'b011001111011101011: begin rgb_reg = 3'b111; end
            18'b011001111011101100: begin rgb_reg = 3'b111; end
            18'b011001111011110100: begin rgb_reg = 3'b111; end
            18'b011001111011110101: begin rgb_reg = 3'b111; end
            18'b011001111011111011: begin rgb_reg = 3'b111; end
            18'b011001111011111100: begin rgb_reg = 3'b111; end
            18'b011001111011111101: begin rgb_reg = 3'b111; end
            18'b011001111011111110: begin rgb_reg = 3'b111; end
            18'b011001111100000010: begin rgb_reg = 3'b111; end
            18'b011001111100000011: begin rgb_reg = 3'b111; end
            18'b011001111100000100: begin rgb_reg = 3'b111; end
            18'b011001111100010001: begin rgb_reg = 3'b111; end
            18'b011001111100010010: begin rgb_reg = 3'b111; end
            18'b011001111100010011: begin rgb_reg = 3'b111; end
            18'b011001111100010100: begin rgb_reg = 3'b111; end
            18'b011001111100010101: begin rgb_reg = 3'b111; end
            18'b011001111100011100: begin rgb_reg = 3'b111; end
            18'b011001111100011101: begin rgb_reg = 3'b111; end
            18'b011001111100011110: begin rgb_reg = 3'b111; end
            18'b011001111100100011: begin rgb_reg = 3'b111; end
            18'b011001111100100100: begin rgb_reg = 3'b111; end
            18'b011001111100100101: begin rgb_reg = 3'b111; end
            18'b011001111100100110: begin rgb_reg = 3'b111; end
            18'b011001111100100111: begin rgb_reg = 3'b111; end
            18'b011001111100101010: begin rgb_reg = 3'b111; end
            18'b011001111100101011: begin rgb_reg = 3'b111; end
            18'b011001111100110011: begin rgb_reg = 3'b111; end
            18'b011001111100110100: begin rgb_reg = 3'b111; end
            18'b011001111100111010: begin rgb_reg = 3'b111; end
            18'b011001111100111011: begin rgb_reg = 3'b111; end
            18'b011001111100111100: begin rgb_reg = 3'b111; end
            18'b011001111100111101: begin rgb_reg = 3'b111; end
            18'b011010000010111110: begin rgb_reg = 3'b111; end
            18'b011010000010111111: begin rgb_reg = 3'b111; end
            18'b011010000011001011: begin rgb_reg = 3'b111; end
            18'b011010000011001100: begin rgb_reg = 3'b111; end
            18'b011010000011001101: begin rgb_reg = 3'b111; end
            18'b011010000011010010: begin rgb_reg = 3'b111; end
            18'b011010000011010011: begin rgb_reg = 3'b111; end
            18'b011010000011010100: begin rgb_reg = 3'b111; end
            18'b011010000011010101: begin rgb_reg = 3'b111; end
            18'b011010000011010110: begin rgb_reg = 3'b111; end
            18'b011010000011100010: begin rgb_reg = 3'b111; end
            18'b011010000011100011: begin rgb_reg = 3'b111; end
            18'b011010000011101011: begin rgb_reg = 3'b111; end
            18'b011010000011101100: begin rgb_reg = 3'b111; end
            18'b011010000011110100: begin rgb_reg = 3'b111; end
            18'b011010000011110101: begin rgb_reg = 3'b111; end
            18'b011010000011111010: begin rgb_reg = 3'b111; end
            18'b011010000011111011: begin rgb_reg = 3'b111; end
            18'b011010000011111100: begin rgb_reg = 3'b111; end
            18'b011010000011111101: begin rgb_reg = 3'b111; end
            18'b011010000011111110: begin rgb_reg = 3'b111; end
            18'b011010000100000001: begin rgb_reg = 3'b111; end
            18'b011010000100000010: begin rgb_reg = 3'b111; end
            18'b011010000100000011: begin rgb_reg = 3'b111; end
            18'b011010000100010011: begin rgb_reg = 3'b111; end
            18'b011010000100010100: begin rgb_reg = 3'b111; end
            18'b011010000100010101: begin rgb_reg = 3'b111; end
            18'b011010000100011100: begin rgb_reg = 3'b111; end
            18'b011010000100011101: begin rgb_reg = 3'b111; end
            18'b011010000100011110: begin rgb_reg = 3'b111; end
            18'b011010000100100011: begin rgb_reg = 3'b111; end
            18'b011010000100100100: begin rgb_reg = 3'b111; end
            18'b011010000100100101: begin rgb_reg = 3'b111; end
            18'b011010000100100110: begin rgb_reg = 3'b111; end
            18'b011010000100100111: begin rgb_reg = 3'b111; end
            18'b011010000100110011: begin rgb_reg = 3'b111; end
            18'b011010000100110100: begin rgb_reg = 3'b111; end
            18'b011010000100111100: begin rgb_reg = 3'b111; end
            18'b011010000100111101: begin rgb_reg = 3'b111; end
            18'b011010001010111110: begin rgb_reg = 3'b111; end
            18'b011010001010111111: begin rgb_reg = 3'b111; end
            18'b011010001011001011: begin rgb_reg = 3'b111; end
            18'b011010001011001100: begin rgb_reg = 3'b111; end
            18'b011010001011001101: begin rgb_reg = 3'b111; end
            18'b011010001011010010: begin rgb_reg = 3'b111; end
            18'b011010001011010011: begin rgb_reg = 3'b111; end
            18'b011010001011010100: begin rgb_reg = 3'b111; end
            18'b011010001011010101: begin rgb_reg = 3'b111; end
            18'b011010001011010110: begin rgb_reg = 3'b111; end
            18'b011010001011100010: begin rgb_reg = 3'b111; end
            18'b011010001011100011: begin rgb_reg = 3'b111; end
            18'b011010001011101011: begin rgb_reg = 3'b111; end
            18'b011010001011101100: begin rgb_reg = 3'b111; end
            18'b011010001011110100: begin rgb_reg = 3'b111; end
            18'b011010001011110101: begin rgb_reg = 3'b111; end
            18'b011010001011111010: begin rgb_reg = 3'b111; end
            18'b011010001011111011: begin rgb_reg = 3'b111; end
            18'b011010001011111100: begin rgb_reg = 3'b111; end
            18'b011010001011111101: begin rgb_reg = 3'b111; end
            18'b011010001011111110: begin rgb_reg = 3'b111; end
            18'b011010001100000001: begin rgb_reg = 3'b111; end
            18'b011010001100000010: begin rgb_reg = 3'b111; end
            18'b011010001100000011: begin rgb_reg = 3'b111; end
            18'b011010001100010011: begin rgb_reg = 3'b111; end
            18'b011010001100010100: begin rgb_reg = 3'b111; end
            18'b011010001100010101: begin rgb_reg = 3'b111; end
            18'b011010001100011100: begin rgb_reg = 3'b111; end
            18'b011010001100011101: begin rgb_reg = 3'b111; end
            18'b011010001100011110: begin rgb_reg = 3'b111; end
            18'b011010001100100011: begin rgb_reg = 3'b111; end
            18'b011010001100100100: begin rgb_reg = 3'b111; end
            18'b011010001100100101: begin rgb_reg = 3'b111; end
            18'b011010001100100110: begin rgb_reg = 3'b111; end
            18'b011010001100100111: begin rgb_reg = 3'b111; end
            18'b011010001100110011: begin rgb_reg = 3'b111; end
            18'b011010001100110100: begin rgb_reg = 3'b111; end
            18'b011010001100111100: begin rgb_reg = 3'b111; end
            18'b011010001100111101: begin rgb_reg = 3'b111; end
            18'b011010010010111110: begin rgb_reg = 3'b111; end
            18'b011010010010111111: begin rgb_reg = 3'b111; end
            18'b011010010011000000: begin rgb_reg = 3'b111; end
            18'b011010010011000001: begin rgb_reg = 3'b111; end
            18'b011010010011000010: begin rgb_reg = 3'b111; end
            18'b011010010011000011: begin rgb_reg = 3'b111; end
            18'b011010010011000100: begin rgb_reg = 3'b111; end
            18'b011010010011000101: begin rgb_reg = 3'b111; end
            18'b011010010011000110: begin rgb_reg = 3'b111; end
            18'b011010010011001011: begin rgb_reg = 3'b111; end
            18'b011010010011001100: begin rgb_reg = 3'b111; end
            18'b011010010011001101: begin rgb_reg = 3'b111; end
            18'b011010010011010000: begin rgb_reg = 3'b111; end
            18'b011010010011010001: begin rgb_reg = 3'b111; end
            18'b011010010011010100: begin rgb_reg = 3'b111; end
            18'b011010010011010101: begin rgb_reg = 3'b111; end
            18'b011010010011010110: begin rgb_reg = 3'b111; end
            18'b011010010011011101: begin rgb_reg = 3'b111; end
            18'b011010010011011110: begin rgb_reg = 3'b111; end
            18'b011010010011011111: begin rgb_reg = 3'b111; end
            18'b011010010011100000: begin rgb_reg = 3'b111; end
            18'b011010010011100001: begin rgb_reg = 3'b111; end
            18'b011010010011101011: begin rgb_reg = 3'b111; end
            18'b011010010011101100: begin rgb_reg = 3'b111; end
            18'b011010010011110100: begin rgb_reg = 3'b111; end
            18'b011010010011110101: begin rgb_reg = 3'b111; end
            18'b011010010011111000: begin rgb_reg = 3'b111; end
            18'b011010010011111001: begin rgb_reg = 3'b111; end
            18'b011010010011111010: begin rgb_reg = 3'b111; end
            18'b011010010011111101: begin rgb_reg = 3'b111; end
            18'b011010010011111110: begin rgb_reg = 3'b111; end
            18'b011010010100000001: begin rgb_reg = 3'b111; end
            18'b011010010100000010: begin rgb_reg = 3'b111; end
            18'b011010010100000011: begin rgb_reg = 3'b111; end
            18'b011010010100000100: begin rgb_reg = 3'b111; end
            18'b011010010100000101: begin rgb_reg = 3'b111; end
            18'b011010010100000110: begin rgb_reg = 3'b111; end
            18'b011010010100000111: begin rgb_reg = 3'b111; end
            18'b011010010100001000: begin rgb_reg = 3'b111; end
            18'b011010010100001001: begin rgb_reg = 3'b111; end
            18'b011010010100010011: begin rgb_reg = 3'b111; end
            18'b011010010100010100: begin rgb_reg = 3'b111; end
            18'b011010010100010101: begin rgb_reg = 3'b111; end
            18'b011010010100011100: begin rgb_reg = 3'b111; end
            18'b011010010100011101: begin rgb_reg = 3'b111; end
            18'b011010010100011110: begin rgb_reg = 3'b111; end
            18'b011010010100100001: begin rgb_reg = 3'b111; end
            18'b011010010100100010: begin rgb_reg = 3'b111; end
            18'b011010010100100101: begin rgb_reg = 3'b111; end
            18'b011010010100100110: begin rgb_reg = 3'b111; end
            18'b011010010100100111: begin rgb_reg = 3'b111; end
            18'b011010010100101110: begin rgb_reg = 3'b111; end
            18'b011010010100101111: begin rgb_reg = 3'b111; end
            18'b011010010100110000: begin rgb_reg = 3'b111; end
            18'b011010010100110001: begin rgb_reg = 3'b111; end
            18'b011010010100110010: begin rgb_reg = 3'b111; end
            18'b011010010100111100: begin rgb_reg = 3'b111; end
            18'b011010010100111101: begin rgb_reg = 3'b111; end
            18'b011010011010111110: begin rgb_reg = 3'b111; end
            18'b011010011010111111: begin rgb_reg = 3'b111; end
            18'b011010011011000000: begin rgb_reg = 3'b111; end
            18'b011010011011000001: begin rgb_reg = 3'b111; end
            18'b011010011011000010: begin rgb_reg = 3'b111; end
            18'b011010011011000011: begin rgb_reg = 3'b111; end
            18'b011010011011000100: begin rgb_reg = 3'b111; end
            18'b011010011011000101: begin rgb_reg = 3'b111; end
            18'b011010011011000110: begin rgb_reg = 3'b111; end
            18'b011010011011001011: begin rgb_reg = 3'b111; end
            18'b011010011011001100: begin rgb_reg = 3'b111; end
            18'b011010011011001101: begin rgb_reg = 3'b111; end
            18'b011010011011010000: begin rgb_reg = 3'b111; end
            18'b011010011011010001: begin rgb_reg = 3'b111; end
            18'b011010011011010100: begin rgb_reg = 3'b111; end
            18'b011010011011010101: begin rgb_reg = 3'b111; end
            18'b011010011011010110: begin rgb_reg = 3'b111; end
            18'b011010011011011101: begin rgb_reg = 3'b111; end
            18'b011010011011011110: begin rgb_reg = 3'b111; end
            18'b011010011011011111: begin rgb_reg = 3'b111; end
            18'b011010011011100000: begin rgb_reg = 3'b111; end
            18'b011010011011100001: begin rgb_reg = 3'b111; end
            18'b011010011011101011: begin rgb_reg = 3'b111; end
            18'b011010011011101100: begin rgb_reg = 3'b111; end
            18'b011010011011110100: begin rgb_reg = 3'b111; end
            18'b011010011011110101: begin rgb_reg = 3'b111; end
            18'b011010011011111000: begin rgb_reg = 3'b111; end
            18'b011010011011111001: begin rgb_reg = 3'b111; end
            18'b011010011011111010: begin rgb_reg = 3'b111; end
            18'b011010011011111101: begin rgb_reg = 3'b111; end
            18'b011010011011111110: begin rgb_reg = 3'b111; end
            18'b011010011100000001: begin rgb_reg = 3'b111; end
            18'b011010011100000010: begin rgb_reg = 3'b111; end
            18'b011010011100000011: begin rgb_reg = 3'b111; end
            18'b011010011100000100: begin rgb_reg = 3'b111; end
            18'b011010011100000101: begin rgb_reg = 3'b111; end
            18'b011010011100000110: begin rgb_reg = 3'b111; end
            18'b011010011100000111: begin rgb_reg = 3'b111; end
            18'b011010011100001000: begin rgb_reg = 3'b111; end
            18'b011010011100001001: begin rgb_reg = 3'b111; end
            18'b011010011100010011: begin rgb_reg = 3'b111; end
            18'b011010011100010100: begin rgb_reg = 3'b111; end
            18'b011010011100010101: begin rgb_reg = 3'b111; end
            18'b011010011100011100: begin rgb_reg = 3'b111; end
            18'b011010011100011101: begin rgb_reg = 3'b111; end
            18'b011010011100011110: begin rgb_reg = 3'b111; end
            18'b011010011100100001: begin rgb_reg = 3'b111; end
            18'b011010011100100010: begin rgb_reg = 3'b111; end
            18'b011010011100100101: begin rgb_reg = 3'b111; end
            18'b011010011100100110: begin rgb_reg = 3'b111; end
            18'b011010011100100111: begin rgb_reg = 3'b111; end
            18'b011010011100101110: begin rgb_reg = 3'b111; end
            18'b011010011100101111: begin rgb_reg = 3'b111; end
            18'b011010011100110000: begin rgb_reg = 3'b111; end
            18'b011010011100110001: begin rgb_reg = 3'b111; end
            18'b011010011100110010: begin rgb_reg = 3'b111; end
            18'b011010011100111100: begin rgb_reg = 3'b111; end
            18'b011010011100111101: begin rgb_reg = 3'b111; end
            18'b011010100010111110: begin rgb_reg = 3'b111; end
            18'b011010100010111111: begin rgb_reg = 3'b111; end
            18'b011010100011000111: begin rgb_reg = 3'b111; end
            18'b011010100011001000: begin rgb_reg = 3'b111; end
            18'b011010100011001011: begin rgb_reg = 3'b111; end
            18'b011010100011001100: begin rgb_reg = 3'b111; end
            18'b011010100011001101: begin rgb_reg = 3'b111; end
            18'b011010100011001110: begin rgb_reg = 3'b111; end
            18'b011010100011001111: begin rgb_reg = 3'b111; end
            18'b011010100011010100: begin rgb_reg = 3'b111; end
            18'b011010100011010101: begin rgb_reg = 3'b111; end
            18'b011010100011010110: begin rgb_reg = 3'b111; end
            18'b011010100011100010: begin rgb_reg = 3'b111; end
            18'b011010100011100011: begin rgb_reg = 3'b111; end
            18'b011010100011101011: begin rgb_reg = 3'b111; end
            18'b011010100011101100: begin rgb_reg = 3'b111; end
            18'b011010100011110100: begin rgb_reg = 3'b111; end
            18'b011010100011110101: begin rgb_reg = 3'b111; end
            18'b011010100011110110: begin rgb_reg = 3'b111; end
            18'b011010100011110111: begin rgb_reg = 3'b111; end
            18'b011010100011111101: begin rgb_reg = 3'b111; end
            18'b011010100011111110: begin rgb_reg = 3'b111; end
            18'b011010100100000001: begin rgb_reg = 3'b111; end
            18'b011010100100000010: begin rgb_reg = 3'b111; end
            18'b011010100100000011: begin rgb_reg = 3'b111; end
            18'b011010100100001010: begin rgb_reg = 3'b111; end
            18'b011010100100001011: begin rgb_reg = 3'b111; end
            18'b011010100100001100: begin rgb_reg = 3'b111; end
            18'b011010100100010011: begin rgb_reg = 3'b111; end
            18'b011010100100010100: begin rgb_reg = 3'b111; end
            18'b011010100100010101: begin rgb_reg = 3'b111; end
            18'b011010100100011100: begin rgb_reg = 3'b111; end
            18'b011010100100011101: begin rgb_reg = 3'b111; end
            18'b011010100100011110: begin rgb_reg = 3'b111; end
            18'b011010100100011111: begin rgb_reg = 3'b111; end
            18'b011010100100100000: begin rgb_reg = 3'b111; end
            18'b011010100100100101: begin rgb_reg = 3'b111; end
            18'b011010100100100110: begin rgb_reg = 3'b111; end
            18'b011010100100100111: begin rgb_reg = 3'b111; end
            18'b011010100100101100: begin rgb_reg = 3'b111; end
            18'b011010100100101101: begin rgb_reg = 3'b111; end
            18'b011010100100111100: begin rgb_reg = 3'b111; end
            18'b011010100100111101: begin rgb_reg = 3'b111; end
            18'b011010101010111110: begin rgb_reg = 3'b111; end
            18'b011010101010111111: begin rgb_reg = 3'b111; end
            18'b011010101011000111: begin rgb_reg = 3'b111; end
            18'b011010101011001000: begin rgb_reg = 3'b111; end
            18'b011010101011001011: begin rgb_reg = 3'b111; end
            18'b011010101011001100: begin rgb_reg = 3'b111; end
            18'b011010101011001101: begin rgb_reg = 3'b111; end
            18'b011010101011001110: begin rgb_reg = 3'b111; end
            18'b011010101011001111: begin rgb_reg = 3'b111; end
            18'b011010101011010100: begin rgb_reg = 3'b111; end
            18'b011010101011010101: begin rgb_reg = 3'b111; end
            18'b011010101011010110: begin rgb_reg = 3'b111; end
            18'b011010101011100010: begin rgb_reg = 3'b111; end
            18'b011010101011100011: begin rgb_reg = 3'b111; end
            18'b011010101011101011: begin rgb_reg = 3'b111; end
            18'b011010101011101100: begin rgb_reg = 3'b111; end
            18'b011010101011110100: begin rgb_reg = 3'b111; end
            18'b011010101011110101: begin rgb_reg = 3'b111; end
            18'b011010101011110110: begin rgb_reg = 3'b111; end
            18'b011010101011110111: begin rgb_reg = 3'b111; end
            18'b011010101011111101: begin rgb_reg = 3'b111; end
            18'b011010101011111110: begin rgb_reg = 3'b111; end
            18'b011010101100000001: begin rgb_reg = 3'b111; end
            18'b011010101100000010: begin rgb_reg = 3'b111; end
            18'b011010101100000011: begin rgb_reg = 3'b111; end
            18'b011010101100001010: begin rgb_reg = 3'b111; end
            18'b011010101100001011: begin rgb_reg = 3'b111; end
            18'b011010101100001100: begin rgb_reg = 3'b111; end
            18'b011010101100010011: begin rgb_reg = 3'b111; end
            18'b011010101100010100: begin rgb_reg = 3'b111; end
            18'b011010101100010101: begin rgb_reg = 3'b111; end
            18'b011010101100011100: begin rgb_reg = 3'b111; end
            18'b011010101100011101: begin rgb_reg = 3'b111; end
            18'b011010101100011110: begin rgb_reg = 3'b111; end
            18'b011010101100011111: begin rgb_reg = 3'b111; end
            18'b011010101100100000: begin rgb_reg = 3'b111; end
            18'b011010101100100101: begin rgb_reg = 3'b111; end
            18'b011010101100100110: begin rgb_reg = 3'b111; end
            18'b011010101100100111: begin rgb_reg = 3'b111; end
            18'b011010101100101100: begin rgb_reg = 3'b111; end
            18'b011010101100101101: begin rgb_reg = 3'b111; end
            18'b011010101100111100: begin rgb_reg = 3'b111; end
            18'b011010101100111101: begin rgb_reg = 3'b111; end
            18'b011010110010111110: begin rgb_reg = 3'b111; end
            18'b011010110010111111: begin rgb_reg = 3'b111; end
            18'b011010110011000111: begin rgb_reg = 3'b111; end
            18'b011010110011001000: begin rgb_reg = 3'b111; end
            18'b011010110011001011: begin rgb_reg = 3'b111; end
            18'b011010110011001100: begin rgb_reg = 3'b111; end
            18'b011010110011001101: begin rgb_reg = 3'b111; end
            18'b011010110011010100: begin rgb_reg = 3'b111; end
            18'b011010110011010101: begin rgb_reg = 3'b111; end
            18'b011010110011010110: begin rgb_reg = 3'b111; end
            18'b011010110011011001: begin rgb_reg = 3'b111; end
            18'b011010110011011010: begin rgb_reg = 3'b111; end
            18'b011010110011100010: begin rgb_reg = 3'b111; end
            18'b011010110011100011: begin rgb_reg = 3'b111; end
            18'b011010110011101011: begin rgb_reg = 3'b111; end
            18'b011010110011101100: begin rgb_reg = 3'b111; end
            18'b011010110011110100: begin rgb_reg = 3'b111; end
            18'b011010110011110101: begin rgb_reg = 3'b111; end
            18'b011010110011111101: begin rgb_reg = 3'b111; end
            18'b011010110011111110: begin rgb_reg = 3'b111; end
            18'b011010110100000001: begin rgb_reg = 3'b111; end
            18'b011010110100000010: begin rgb_reg = 3'b111; end
            18'b011010110100000011: begin rgb_reg = 3'b111; end
            18'b011010110100001010: begin rgb_reg = 3'b111; end
            18'b011010110100001011: begin rgb_reg = 3'b111; end
            18'b011010110100001100: begin rgb_reg = 3'b111; end
            18'b011010110100010011: begin rgb_reg = 3'b111; end
            18'b011010110100010100: begin rgb_reg = 3'b111; end
            18'b011010110100010101: begin rgb_reg = 3'b111; end
            18'b011010110100011100: begin rgb_reg = 3'b111; end
            18'b011010110100011101: begin rgb_reg = 3'b111; end
            18'b011010110100011110: begin rgb_reg = 3'b111; end
            18'b011010110100100101: begin rgb_reg = 3'b111; end
            18'b011010110100100110: begin rgb_reg = 3'b111; end
            18'b011010110100100111: begin rgb_reg = 3'b111; end
            18'b011010110100101010: begin rgb_reg = 3'b111; end
            18'b011010110100101011: begin rgb_reg = 3'b111; end
            18'b011010110100111100: begin rgb_reg = 3'b111; end
            18'b011010110100111101: begin rgb_reg = 3'b111; end
            18'b011010111010111110: begin rgb_reg = 3'b111; end
            18'b011010111010111111: begin rgb_reg = 3'b111; end
            18'b011010111011000111: begin rgb_reg = 3'b111; end
            18'b011010111011001000: begin rgb_reg = 3'b111; end
            18'b011010111011001011: begin rgb_reg = 3'b111; end
            18'b011010111011001100: begin rgb_reg = 3'b111; end
            18'b011010111011001101: begin rgb_reg = 3'b111; end
            18'b011010111011010100: begin rgb_reg = 3'b111; end
            18'b011010111011010101: begin rgb_reg = 3'b111; end
            18'b011010111011010110: begin rgb_reg = 3'b111; end
            18'b011010111011011001: begin rgb_reg = 3'b111; end
            18'b011010111011011010: begin rgb_reg = 3'b111; end
            18'b011010111011100010: begin rgb_reg = 3'b111; end
            18'b011010111011100011: begin rgb_reg = 3'b111; end
            18'b011010111011101011: begin rgb_reg = 3'b111; end
            18'b011010111011101100: begin rgb_reg = 3'b111; end
            18'b011010111011110100: begin rgb_reg = 3'b111; end
            18'b011010111011110101: begin rgb_reg = 3'b111; end
            18'b011010111011111101: begin rgb_reg = 3'b111; end
            18'b011010111011111110: begin rgb_reg = 3'b111; end
            18'b011010111100000001: begin rgb_reg = 3'b111; end
            18'b011010111100000010: begin rgb_reg = 3'b111; end
            18'b011010111100000011: begin rgb_reg = 3'b111; end
            18'b011010111100001010: begin rgb_reg = 3'b111; end
            18'b011010111100001011: begin rgb_reg = 3'b111; end
            18'b011010111100001100: begin rgb_reg = 3'b111; end
            18'b011010111100010011: begin rgb_reg = 3'b111; end
            18'b011010111100010100: begin rgb_reg = 3'b111; end
            18'b011010111100010101: begin rgb_reg = 3'b111; end
            18'b011010111100011100: begin rgb_reg = 3'b111; end
            18'b011010111100011101: begin rgb_reg = 3'b111; end
            18'b011010111100011110: begin rgb_reg = 3'b111; end
            18'b011010111100100101: begin rgb_reg = 3'b111; end
            18'b011010111100100110: begin rgb_reg = 3'b111; end
            18'b011010111100100111: begin rgb_reg = 3'b111; end
            18'b011010111100101010: begin rgb_reg = 3'b111; end
            18'b011010111100101011: begin rgb_reg = 3'b111; end
            18'b011010111100111100: begin rgb_reg = 3'b111; end
            18'b011010111100111101: begin rgb_reg = 3'b111; end
            18'b011011000010111110: begin rgb_reg = 3'b111; end
            18'b011011000010111111: begin rgb_reg = 3'b111; end
            18'b011011000011000000: begin rgb_reg = 3'b111; end
            18'b011011000011000001: begin rgb_reg = 3'b111; end
            18'b011011000011000010: begin rgb_reg = 3'b111; end
            18'b011011000011000011: begin rgb_reg = 3'b111; end
            18'b011011000011000100: begin rgb_reg = 3'b111; end
            18'b011011000011000101: begin rgb_reg = 3'b111; end
            18'b011011000011000110: begin rgb_reg = 3'b111; end
            18'b011011000011000111: begin rgb_reg = 3'b111; end
            18'b011011000011001000: begin rgb_reg = 3'b111; end
            18'b011011000011001100: begin rgb_reg = 3'b111; end
            18'b011011000011001101: begin rgb_reg = 3'b111; end
            18'b011011000011001110: begin rgb_reg = 3'b111; end
            18'b011011000011001111: begin rgb_reg = 3'b111; end
            18'b011011000011010000: begin rgb_reg = 3'b111; end
            18'b011011000011010001: begin rgb_reg = 3'b111; end
            18'b011011000011010010: begin rgb_reg = 3'b111; end
            18'b011011000011010011: begin rgb_reg = 3'b111; end
            18'b011011000011010100: begin rgb_reg = 3'b111; end
            18'b011011000011010101: begin rgb_reg = 3'b111; end
            18'b011011000011011001: begin rgb_reg = 3'b111; end
            18'b011011000011011010: begin rgb_reg = 3'b111; end
            18'b011011000011011011: begin rgb_reg = 3'b111; end
            18'b011011000011011100: begin rgb_reg = 3'b111; end
            18'b011011000011011101: begin rgb_reg = 3'b111; end
            18'b011011000011011110: begin rgb_reg = 3'b111; end
            18'b011011000011011111: begin rgb_reg = 3'b111; end
            18'b011011000011100000: begin rgb_reg = 3'b111; end
            18'b011011000011100001: begin rgb_reg = 3'b111; end
            18'b011011000011100010: begin rgb_reg = 3'b111; end
            18'b011011000011100011: begin rgb_reg = 3'b111; end
            18'b011011000011100111: begin rgb_reg = 3'b111; end
            18'b011011000011101000: begin rgb_reg = 3'b111; end
            18'b011011000011101001: begin rgb_reg = 3'b111; end
            18'b011011000011101010: begin rgb_reg = 3'b111; end
            18'b011011000011101011: begin rgb_reg = 3'b111; end
            18'b011011000011101100: begin rgb_reg = 3'b111; end
            18'b011011000011101101: begin rgb_reg = 3'b111; end
            18'b011011000011101110: begin rgb_reg = 3'b111; end
            18'b011011000011101111: begin rgb_reg = 3'b111; end
            18'b011011000011110000: begin rgb_reg = 3'b111; end
            18'b011011000011110100: begin rgb_reg = 3'b111; end
            18'b011011000011110101: begin rgb_reg = 3'b111; end
            18'b011011000011110110: begin rgb_reg = 3'b111; end
            18'b011011000011110111: begin rgb_reg = 3'b111; end
            18'b011011000011111000: begin rgb_reg = 3'b111; end
            18'b011011000011111001: begin rgb_reg = 3'b111; end
            18'b011011000011111010: begin rgb_reg = 3'b111; end
            18'b011011000011111011: begin rgb_reg = 3'b111; end
            18'b011011000011111100: begin rgb_reg = 3'b111; end
            18'b011011000011111101: begin rgb_reg = 3'b111; end
            18'b011011000011111110: begin rgb_reg = 3'b111; end
            18'b011011000100000010: begin rgb_reg = 3'b111; end
            18'b011011000100000011: begin rgb_reg = 3'b111; end
            18'b011011000100000100: begin rgb_reg = 3'b111; end
            18'b011011000100000101: begin rgb_reg = 3'b111; end
            18'b011011000100000110: begin rgb_reg = 3'b111; end
            18'b011011000100000111: begin rgb_reg = 3'b111; end
            18'b011011000100001000: begin rgb_reg = 3'b111; end
            18'b011011000100001001: begin rgb_reg = 3'b111; end
            18'b011011000100001010: begin rgb_reg = 3'b111; end
            18'b011011000100001011: begin rgb_reg = 3'b111; end
            18'b011011000100001111: begin rgb_reg = 3'b111; end
            18'b011011000100010000: begin rgb_reg = 3'b111; end
            18'b011011000100010001: begin rgb_reg = 3'b111; end
            18'b011011000100010010: begin rgb_reg = 3'b111; end
            18'b011011000100010011: begin rgb_reg = 3'b111; end
            18'b011011000100010100: begin rgb_reg = 3'b111; end
            18'b011011000100010101: begin rgb_reg = 3'b111; end
            18'b011011000100010110: begin rgb_reg = 3'b111; end
            18'b011011000100010111: begin rgb_reg = 3'b111; end
            18'b011011000100011000: begin rgb_reg = 3'b111; end
            18'b011011000100011001: begin rgb_reg = 3'b111; end
            18'b011011000100011101: begin rgb_reg = 3'b111; end
            18'b011011000100011110: begin rgb_reg = 3'b111; end
            18'b011011000100011111: begin rgb_reg = 3'b111; end
            18'b011011000100100000: begin rgb_reg = 3'b111; end
            18'b011011000100100001: begin rgb_reg = 3'b111; end
            18'b011011000100100010: begin rgb_reg = 3'b111; end
            18'b011011000100100011: begin rgb_reg = 3'b111; end
            18'b011011000100100100: begin rgb_reg = 3'b111; end
            18'b011011000100100101: begin rgb_reg = 3'b111; end
            18'b011011000100100110: begin rgb_reg = 3'b111; end
            18'b011011000100101010: begin rgb_reg = 3'b111; end
            18'b011011000100101011: begin rgb_reg = 3'b111; end
            18'b011011000100101100: begin rgb_reg = 3'b111; end
            18'b011011000100101101: begin rgb_reg = 3'b111; end
            18'b011011000100101110: begin rgb_reg = 3'b111; end
            18'b011011000100101111: begin rgb_reg = 3'b111; end
            18'b011011000100110000: begin rgb_reg = 3'b111; end
            18'b011011000100110001: begin rgb_reg = 3'b111; end
            18'b011011000100110010: begin rgb_reg = 3'b111; end
            18'b011011000100110011: begin rgb_reg = 3'b111; end
            18'b011011000100110100: begin rgb_reg = 3'b111; end
            18'b011011000100111000: begin rgb_reg = 3'b111; end
            18'b011011000100111001: begin rgb_reg = 3'b111; end
            18'b011011000100111010: begin rgb_reg = 3'b111; end
            18'b011011000100111011: begin rgb_reg = 3'b111; end
            18'b011011000100111100: begin rgb_reg = 3'b111; end
            18'b011011000100111101: begin rgb_reg = 3'b111; end
            18'b011011000100111110: begin rgb_reg = 3'b111; end
            18'b011011000100111111: begin rgb_reg = 3'b111; end
            18'b011011000101000000: begin rgb_reg = 3'b111; end
            18'b011011000101000001: begin rgb_reg = 3'b111; end
            18'b011011001011000000: begin rgb_reg = 3'b111; end
            18'b011011001011000001: begin rgb_reg = 3'b111; end
            18'b011011001011000010: begin rgb_reg = 3'b111; end
            18'b011011001011000011: begin rgb_reg = 3'b111; end
            18'b011011001011000100: begin rgb_reg = 3'b111; end
            18'b011011001011000101: begin rgb_reg = 3'b111; end
            18'b011011001011000110: begin rgb_reg = 3'b111; end
            18'b011011001011001101: begin rgb_reg = 3'b111; end
            18'b011011001011001110: begin rgb_reg = 3'b111; end
            18'b011011001011001111: begin rgb_reg = 3'b111; end
            18'b011011001011010000: begin rgb_reg = 3'b111; end
            18'b011011001011010001: begin rgb_reg = 3'b111; end
            18'b011011001011010010: begin rgb_reg = 3'b111; end
            18'b011011001011010011: begin rgb_reg = 3'b111; end
            18'b011011001011011011: begin rgb_reg = 3'b111; end
            18'b011011001011011100: begin rgb_reg = 3'b111; end
            18'b011011001011011101: begin rgb_reg = 3'b111; end
            18'b011011001011011110: begin rgb_reg = 3'b111; end
            18'b011011001011011111: begin rgb_reg = 3'b111; end
            18'b011011001011100000: begin rgb_reg = 3'b111; end
            18'b011011001011100001: begin rgb_reg = 3'b111; end
            18'b011011001011100110: begin rgb_reg = 3'b111; end
            18'b011011001011100111: begin rgb_reg = 3'b111; end
            18'b011011001011101000: begin rgb_reg = 3'b111; end
            18'b011011001011101001: begin rgb_reg = 3'b111; end
            18'b011011001011101010: begin rgb_reg = 3'b111; end
            18'b011011001011101011: begin rgb_reg = 3'b111; end
            18'b011011001011101100: begin rgb_reg = 3'b111; end
            18'b011011001011101101: begin rgb_reg = 3'b111; end
            18'b011011001011101110: begin rgb_reg = 3'b111; end
            18'b011011001011101111: begin rgb_reg = 3'b111; end
            18'b011011001011110000: begin rgb_reg = 3'b111; end
            18'b011011001011110001: begin rgb_reg = 3'b111; end
            18'b011011001011110110: begin rgb_reg = 3'b111; end
            18'b011011001011110111: begin rgb_reg = 3'b111; end
            18'b011011001011111000: begin rgb_reg = 3'b111; end
            18'b011011001011111001: begin rgb_reg = 3'b111; end
            18'b011011001011111010: begin rgb_reg = 3'b111; end
            18'b011011001011111011: begin rgb_reg = 3'b111; end
            18'b011011001011111100: begin rgb_reg = 3'b111; end
            18'b011011001100000011: begin rgb_reg = 3'b111; end
            18'b011011001100000100: begin rgb_reg = 3'b111; end
            18'b011011001100000101: begin rgb_reg = 3'b111; end
            18'b011011001100000110: begin rgb_reg = 3'b111; end
            18'b011011001100000111: begin rgb_reg = 3'b111; end
            18'b011011001100001000: begin rgb_reg = 3'b111; end
            18'b011011001100001001: begin rgb_reg = 3'b111; end
            18'b011011001100001111: begin rgb_reg = 3'b111; end
            18'b011011001100010000: begin rgb_reg = 3'b111; end
            18'b011011001100010001: begin rgb_reg = 3'b111; end
            18'b011011001100010010: begin rgb_reg = 3'b111; end
            18'b011011001100010011: begin rgb_reg = 3'b111; end
            18'b011011001100010100: begin rgb_reg = 3'b111; end
            18'b011011001100010101: begin rgb_reg = 3'b111; end
            18'b011011001100010110: begin rgb_reg = 3'b111; end
            18'b011011001100010111: begin rgb_reg = 3'b111; end
            18'b011011001100011000: begin rgb_reg = 3'b111; end
            18'b011011001100011001: begin rgb_reg = 3'b111; end
            18'b011011001100011110: begin rgb_reg = 3'b111; end
            18'b011011001100011111: begin rgb_reg = 3'b111; end
            18'b011011001100100000: begin rgb_reg = 3'b111; end
            18'b011011001100100001: begin rgb_reg = 3'b111; end
            18'b011011001100100010: begin rgb_reg = 3'b111; end
            18'b011011001100100011: begin rgb_reg = 3'b111; end
            18'b011011001100100100: begin rgb_reg = 3'b111; end
            18'b011011001100101010: begin rgb_reg = 3'b111; end
            18'b011011001100101011: begin rgb_reg = 3'b111; end
            18'b011011001100101100: begin rgb_reg = 3'b111; end
            18'b011011001100101101: begin rgb_reg = 3'b111; end
            18'b011011001100101110: begin rgb_reg = 3'b111; end
            18'b011011001100101111: begin rgb_reg = 3'b111; end
            18'b011011001100110000: begin rgb_reg = 3'b111; end
            18'b011011001100110001: begin rgb_reg = 3'b111; end
            18'b011011001100110010: begin rgb_reg = 3'b111; end
            18'b011011001100110011: begin rgb_reg = 3'b111; end
            18'b011011001100110100: begin rgb_reg = 3'b111; end
            18'b011011001100110111: begin rgb_reg = 3'b111; end
            18'b011011001100111000: begin rgb_reg = 3'b111; end
            18'b011011001100111001: begin rgb_reg = 3'b111; end
            18'b011011001100111010: begin rgb_reg = 3'b111; end
            18'b011011001100111011: begin rgb_reg = 3'b111; end
            18'b011011001100111100: begin rgb_reg = 3'b111; end
            18'b011011001100111101: begin rgb_reg = 3'b111; end
            18'b011011001100111110: begin rgb_reg = 3'b111; end
            18'b011011001100111111: begin rgb_reg = 3'b111; end
            18'b011011001101000000: begin rgb_reg = 3'b111; end
            18'b011011001101000001: begin rgb_reg = 3'b111; end
            18'b011011001101000010: begin rgb_reg = 3'b111; end
            18'b011011010011000000: begin rgb_reg = 3'b111; end
            18'b011011010011000001: begin rgb_reg = 3'b111; end
            18'b011011010011000010: begin rgb_reg = 3'b111; end
            18'b011011010011000011: begin rgb_reg = 3'b111; end
            18'b011011010011000100: begin rgb_reg = 3'b111; end
            18'b011011010011000101: begin rgb_reg = 3'b111; end
            18'b011011010011000110: begin rgb_reg = 3'b111; end
            18'b011011010011001110: begin rgb_reg = 3'b111; end
            18'b011011010011001111: begin rgb_reg = 3'b111; end
            18'b011011010011010000: begin rgb_reg = 3'b111; end
            18'b011011010011010001: begin rgb_reg = 3'b111; end
            18'b011011010011010010: begin rgb_reg = 3'b111; end
            18'b011011010011010011: begin rgb_reg = 3'b111; end
            18'b011011010011011011: begin rgb_reg = 3'b111; end
            18'b011011010011011100: begin rgb_reg = 3'b111; end
            18'b011011010011011101: begin rgb_reg = 3'b111; end
            18'b011011010011011110: begin rgb_reg = 3'b111; end
            18'b011011010011011111: begin rgb_reg = 3'b111; end
            18'b011011010011100000: begin rgb_reg = 3'b111; end
            18'b011011010011100001: begin rgb_reg = 3'b111; end
            18'b011011010011100110: begin rgb_reg = 3'b111; end
            18'b011011010011100111: begin rgb_reg = 3'b111; end
            18'b011011010011101000: begin rgb_reg = 3'b111; end
            18'b011011010011101001: begin rgb_reg = 3'b111; end
            18'b011011010011101010: begin rgb_reg = 3'b111; end
            18'b011011010011101011: begin rgb_reg = 3'b111; end
            18'b011011010011101100: begin rgb_reg = 3'b111; end
            18'b011011010011101101: begin rgb_reg = 3'b111; end
            18'b011011010011101110: begin rgb_reg = 3'b111; end
            18'b011011010011101111: begin rgb_reg = 3'b111; end
            18'b011011010011110000: begin rgb_reg = 3'b111; end
            18'b011011010011110110: begin rgb_reg = 3'b111; end
            18'b011011010011110111: begin rgb_reg = 3'b111; end
            18'b011011010011111000: begin rgb_reg = 3'b111; end
            18'b011011010011111001: begin rgb_reg = 3'b111; end
            18'b011011010011111010: begin rgb_reg = 3'b111; end
            18'b011011010011111011: begin rgb_reg = 3'b111; end
            18'b011011010011111100: begin rgb_reg = 3'b111; end
            18'b011011010100000100: begin rgb_reg = 3'b111; end
            18'b011011010100000101: begin rgb_reg = 3'b111; end
            18'b011011010100000110: begin rgb_reg = 3'b111; end
            18'b011011010100000111: begin rgb_reg = 3'b111; end
            18'b011011010100001000: begin rgb_reg = 3'b111; end
            18'b011011010100001001: begin rgb_reg = 3'b111; end
            18'b011011010100001111: begin rgb_reg = 3'b111; end
            18'b011011010100010000: begin rgb_reg = 3'b111; end
            18'b011011010100010001: begin rgb_reg = 3'b111; end
            18'b011011010100010010: begin rgb_reg = 3'b111; end
            18'b011011010100010011: begin rgb_reg = 3'b111; end
            18'b011011010100010100: begin rgb_reg = 3'b111; end
            18'b011011010100010101: begin rgb_reg = 3'b111; end
            18'b011011010100010110: begin rgb_reg = 3'b111; end
            18'b011011010100010111: begin rgb_reg = 3'b111; end
            18'b011011010100011000: begin rgb_reg = 3'b111; end
            18'b011011010100011001: begin rgb_reg = 3'b111; end
            18'b011011010100011111: begin rgb_reg = 3'b111; end
            18'b011011010100100000: begin rgb_reg = 3'b111; end
            18'b011011010100100001: begin rgb_reg = 3'b111; end
            18'b011011010100100010: begin rgb_reg = 3'b111; end
            18'b011011010100100011: begin rgb_reg = 3'b111; end
            18'b011011010100100100: begin rgb_reg = 3'b111; end
            18'b011011010100101010: begin rgb_reg = 3'b111; end
            18'b011011010100101011: begin rgb_reg = 3'b111; end
            18'b011011010100101100: begin rgb_reg = 3'b111; end
            18'b011011010100101101: begin rgb_reg = 3'b111; end
            18'b011011010100101110: begin rgb_reg = 3'b111; end
            18'b011011010100101111: begin rgb_reg = 3'b111; end
            18'b011011010100110000: begin rgb_reg = 3'b111; end
            18'b011011010100110001: begin rgb_reg = 3'b111; end
            18'b011011010100110010: begin rgb_reg = 3'b111; end
            18'b011011010100110011: begin rgb_reg = 3'b111; end
            18'b011011010100110100: begin rgb_reg = 3'b111; end
            18'b011011010100110111: begin rgb_reg = 3'b111; end
            18'b011011010100111000: begin rgb_reg = 3'b111; end
            18'b011011010100111001: begin rgb_reg = 3'b111; end
            18'b011011010100111010: begin rgb_reg = 3'b111; end
            18'b011011010100111011: begin rgb_reg = 3'b111; end
            18'b011011010100111100: begin rgb_reg = 3'b111; end
            18'b011011010100111101: begin rgb_reg = 3'b111; end
            18'b011011010100111110: begin rgb_reg = 3'b111; end
            18'b011011010100111111: begin rgb_reg = 3'b111; end
            18'b011011010101000000: begin rgb_reg = 3'b111; end
            18'b011011010101000001: begin rgb_reg = 3'b111; end
            18'b011100010010110011: begin rgb_reg = 3'b111; end
            18'b011100010010110100: begin rgb_reg = 3'b111; end
            18'b011100010010110101: begin rgb_reg = 3'b111; end
            18'b011100010010110110: begin rgb_reg = 3'b111; end
            18'b011100010010110111: begin rgb_reg = 3'b111; end
            18'b011100010010111000: begin rgb_reg = 3'b111; end
            18'b011100010011101101: begin rgb_reg = 3'b111; end
            18'b011100010011101110: begin rgb_reg = 3'b111; end
            18'b011100010011110101: begin rgb_reg = 3'b111; end
            18'b011100010011110110: begin rgb_reg = 3'b111; end
            18'b011100010100000111: begin rgb_reg = 3'b111; end
            18'b011100010100001000: begin rgb_reg = 3'b111; end
            18'b011100010100001101: begin rgb_reg = 3'b111; end
            18'b011100010100001110: begin rgb_reg = 3'b111; end
            18'b011100010100111111: begin rgb_reg = 3'b111; end
            18'b011100010101000000: begin rgb_reg = 3'b111; end
            18'b011100011010110011: begin rgb_reg = 3'b111; end
            18'b011100011010110100: begin rgb_reg = 3'b111; end
            18'b011100011010110101: begin rgb_reg = 3'b111; end
            18'b011100011010110110: begin rgb_reg = 3'b111; end
            18'b011100011010110111: begin rgb_reg = 3'b111; end
            18'b011100011010111000: begin rgb_reg = 3'b111; end
            18'b011100011011101101: begin rgb_reg = 3'b111; end
            18'b011100011011101110: begin rgb_reg = 3'b111; end
            18'b011100011011110101: begin rgb_reg = 3'b111; end
            18'b011100011011110110: begin rgb_reg = 3'b111; end
            18'b011100011100000111: begin rgb_reg = 3'b111; end
            18'b011100011100001000: begin rgb_reg = 3'b111; end
            18'b011100011100001101: begin rgb_reg = 3'b111; end
            18'b011100011100001110: begin rgb_reg = 3'b111; end
            18'b011100011100111111: begin rgb_reg = 3'b111; end
            18'b011100011101000000: begin rgb_reg = 3'b111; end
            18'b011100100010110001: begin rgb_reg = 3'b111; end
            18'b011100100010110010: begin rgb_reg = 3'b111; end
            18'b011100100010111001: begin rgb_reg = 3'b111; end
            18'b011100100010111010: begin rgb_reg = 3'b111; end
            18'b011100100011101101: begin rgb_reg = 3'b111; end
            18'b011100100011101110: begin rgb_reg = 3'b111; end
            18'b011100100011101111: begin rgb_reg = 3'b111; end
            18'b011100100011110000: begin rgb_reg = 3'b111; end
            18'b011100100011110011: begin rgb_reg = 3'b111; end
            18'b011100100011110100: begin rgb_reg = 3'b111; end
            18'b011100100011110101: begin rgb_reg = 3'b111; end
            18'b011100100011110110: begin rgb_reg = 3'b111; end
            18'b011100100100000101: begin rgb_reg = 3'b111; end
            18'b011100100100000110: begin rgb_reg = 3'b111; end
            18'b011100100100000111: begin rgb_reg = 3'b111; end
            18'b011100100100001000: begin rgb_reg = 3'b111; end
            18'b011100100100001001: begin rgb_reg = 3'b111; end
            18'b011100100100001010: begin rgb_reg = 3'b111; end
            18'b011100100100001101: begin rgb_reg = 3'b111; end
            18'b011100100100001110: begin rgb_reg = 3'b111; end
            18'b011100100100111101: begin rgb_reg = 3'b111; end
            18'b011100100100111110: begin rgb_reg = 3'b111; end
            18'b011100100100111111: begin rgb_reg = 3'b111; end
            18'b011100100101000000: begin rgb_reg = 3'b111; end
            18'b011100100101000001: begin rgb_reg = 3'b111; end
            18'b011100100101000010: begin rgb_reg = 3'b111; end
            18'b011100101010110001: begin rgb_reg = 3'b111; end
            18'b011100101010110010: begin rgb_reg = 3'b111; end
            18'b011100101010111001: begin rgb_reg = 3'b111; end
            18'b011100101010111010: begin rgb_reg = 3'b111; end
            18'b011100101011101101: begin rgb_reg = 3'b111; end
            18'b011100101011101110: begin rgb_reg = 3'b111; end
            18'b011100101011101111: begin rgb_reg = 3'b111; end
            18'b011100101011110000: begin rgb_reg = 3'b111; end
            18'b011100101011110011: begin rgb_reg = 3'b111; end
            18'b011100101011110100: begin rgb_reg = 3'b111; end
            18'b011100101011110101: begin rgb_reg = 3'b111; end
            18'b011100101011110110: begin rgb_reg = 3'b111; end
            18'b011100101100000101: begin rgb_reg = 3'b111; end
            18'b011100101100000110: begin rgb_reg = 3'b111; end
            18'b011100101100000111: begin rgb_reg = 3'b111; end
            18'b011100101100001000: begin rgb_reg = 3'b111; end
            18'b011100101100001001: begin rgb_reg = 3'b111; end
            18'b011100101100001010: begin rgb_reg = 3'b111; end
            18'b011100101100001101: begin rgb_reg = 3'b111; end
            18'b011100101100001110: begin rgb_reg = 3'b111; end
            18'b011100101100111101: begin rgb_reg = 3'b111; end
            18'b011100101100111110: begin rgb_reg = 3'b111; end
            18'b011100101100111111: begin rgb_reg = 3'b111; end
            18'b011100101101000000: begin rgb_reg = 3'b111; end
            18'b011100101101000001: begin rgb_reg = 3'b111; end
            18'b011100101101000010: begin rgb_reg = 3'b111; end
            18'b011100110010110001: begin rgb_reg = 3'b111; end
            18'b011100110010110010: begin rgb_reg = 3'b111; end
            18'b011100110010110011: begin rgb_reg = 3'b111; end
            18'b011100110010110100: begin rgb_reg = 3'b111; end
            18'b011100110010110101: begin rgb_reg = 3'b111; end
            18'b011100110010110110: begin rgb_reg = 3'b111; end
            18'b011100110010110111: begin rgb_reg = 3'b111; end
            18'b011100110010111000: begin rgb_reg = 3'b111; end
            18'b011100110010111001: begin rgb_reg = 3'b111; end
            18'b011100110010111010: begin rgb_reg = 3'b111; end
            18'b011100110010111101: begin rgb_reg = 3'b111; end
            18'b011100110010111110: begin rgb_reg = 3'b111; end
            18'b011100110010111111: begin rgb_reg = 3'b111; end
            18'b011100110011000000: begin rgb_reg = 3'b111; end
            18'b011100110011000001: begin rgb_reg = 3'b111; end
            18'b011100110011000010: begin rgb_reg = 3'b111; end
            18'b011100110011000011: begin rgb_reg = 3'b111; end
            18'b011100110011000100: begin rgb_reg = 3'b111; end
            18'b011100110011001011: begin rgb_reg = 3'b111; end
            18'b011100110011001100: begin rgb_reg = 3'b111; end
            18'b011100110011001101: begin rgb_reg = 3'b111; end
            18'b011100110011001110: begin rgb_reg = 3'b111; end
            18'b011100110011001111: begin rgb_reg = 3'b111; end
            18'b011100110011010000: begin rgb_reg = 3'b111; end
            18'b011100110011010101: begin rgb_reg = 3'b111; end
            18'b011100110011010110: begin rgb_reg = 3'b111; end
            18'b011100110011010111: begin rgb_reg = 3'b111; end
            18'b011100110011011000: begin rgb_reg = 3'b111; end
            18'b011100110011011001: begin rgb_reg = 3'b111; end
            18'b011100110011011010: begin rgb_reg = 3'b111; end
            18'b011100110011011011: begin rgb_reg = 3'b111; end
            18'b011100110011011100: begin rgb_reg = 3'b111; end
            18'b011100110011101101: begin rgb_reg = 3'b111; end
            18'b011100110011101110: begin rgb_reg = 3'b111; end
            18'b011100110011110001: begin rgb_reg = 3'b111; end
            18'b011100110011110010: begin rgb_reg = 3'b111; end
            18'b011100110011110101: begin rgb_reg = 3'b111; end
            18'b011100110011110110: begin rgb_reg = 3'b111; end
            18'b011100110011111011: begin rgb_reg = 3'b111; end
            18'b011100110011111100: begin rgb_reg = 3'b111; end
            18'b011100110011111101: begin rgb_reg = 3'b111; end
            18'b011100110011111110: begin rgb_reg = 3'b111; end
            18'b011100110011111111: begin rgb_reg = 3'b111; end
            18'b011100110100000000: begin rgb_reg = 3'b111; end
            18'b011100110100000111: begin rgb_reg = 3'b111; end
            18'b011100110100001000: begin rgb_reg = 3'b111; end
            18'b011100110100001101: begin rgb_reg = 3'b111; end
            18'b011100110100001110: begin rgb_reg = 3'b111; end
            18'b011100110100010001: begin rgb_reg = 3'b111; end
            18'b011100110100010010: begin rgb_reg = 3'b111; end
            18'b011100110100010011: begin rgb_reg = 3'b111; end
            18'b011100110100010100: begin rgb_reg = 3'b111; end
            18'b011100110100011011: begin rgb_reg = 3'b111; end
            18'b011100110100011100: begin rgb_reg = 3'b111; end
            18'b011100110100011101: begin rgb_reg = 3'b111; end
            18'b011100110100011110: begin rgb_reg = 3'b111; end
            18'b011100110100011111: begin rgb_reg = 3'b111; end
            18'b011100110100100000: begin rgb_reg = 3'b111; end
            18'b011100110100100111: begin rgb_reg = 3'b111; end
            18'b011100110100101000: begin rgb_reg = 3'b111; end
            18'b011100110100101001: begin rgb_reg = 3'b111; end
            18'b011100110100101010: begin rgb_reg = 3'b111; end
            18'b011100110100101011: begin rgb_reg = 3'b111; end
            18'b011100110100101100: begin rgb_reg = 3'b111; end
            18'b011100110100101101: begin rgb_reg = 3'b111; end
            18'b011100110100101110: begin rgb_reg = 3'b111; end
            18'b011100110100110011: begin rgb_reg = 3'b111; end
            18'b011100110100110100: begin rgb_reg = 3'b111; end
            18'b011100110100110101: begin rgb_reg = 3'b111; end
            18'b011100110100110110: begin rgb_reg = 3'b111; end
            18'b011100110100110111: begin rgb_reg = 3'b111; end
            18'b011100110100111000: begin rgb_reg = 3'b111; end
            18'b011100110100111111: begin rgb_reg = 3'b111; end
            18'b011100110101000000: begin rgb_reg = 3'b111; end
            18'b011100110101000111: begin rgb_reg = 3'b111; end
            18'b011100110101001000: begin rgb_reg = 3'b111; end
            18'b011100110101001001: begin rgb_reg = 3'b111; end
            18'b011100110101001010: begin rgb_reg = 3'b111; end
            18'b011100110101001011: begin rgb_reg = 3'b111; end
            18'b011100110101001100: begin rgb_reg = 3'b111; end
            18'b011100111010110001: begin rgb_reg = 3'b111; end
            18'b011100111010110010: begin rgb_reg = 3'b111; end
            18'b011100111010110011: begin rgb_reg = 3'b111; end
            18'b011100111010110100: begin rgb_reg = 3'b111; end
            18'b011100111010110101: begin rgb_reg = 3'b111; end
            18'b011100111010110110: begin rgb_reg = 3'b111; end
            18'b011100111010110111: begin rgb_reg = 3'b111; end
            18'b011100111010111000: begin rgb_reg = 3'b111; end
            18'b011100111010111001: begin rgb_reg = 3'b111; end
            18'b011100111010111010: begin rgb_reg = 3'b111; end
            18'b011100111010111101: begin rgb_reg = 3'b111; end
            18'b011100111010111110: begin rgb_reg = 3'b111; end
            18'b011100111010111111: begin rgb_reg = 3'b111; end
            18'b011100111011000000: begin rgb_reg = 3'b111; end
            18'b011100111011000001: begin rgb_reg = 3'b111; end
            18'b011100111011000010: begin rgb_reg = 3'b111; end
            18'b011100111011000011: begin rgb_reg = 3'b111; end
            18'b011100111011000100: begin rgb_reg = 3'b111; end
            18'b011100111011001011: begin rgb_reg = 3'b111; end
            18'b011100111011001100: begin rgb_reg = 3'b111; end
            18'b011100111011001101: begin rgb_reg = 3'b111; end
            18'b011100111011001110: begin rgb_reg = 3'b111; end
            18'b011100111011001111: begin rgb_reg = 3'b111; end
            18'b011100111011010000: begin rgb_reg = 3'b111; end
            18'b011100111011010101: begin rgb_reg = 3'b111; end
            18'b011100111011010110: begin rgb_reg = 3'b111; end
            18'b011100111011010111: begin rgb_reg = 3'b111; end
            18'b011100111011011000: begin rgb_reg = 3'b111; end
            18'b011100111011011001: begin rgb_reg = 3'b111; end
            18'b011100111011011010: begin rgb_reg = 3'b111; end
            18'b011100111011011011: begin rgb_reg = 3'b111; end
            18'b011100111011011100: begin rgb_reg = 3'b111; end
            18'b011100111011101101: begin rgb_reg = 3'b111; end
            18'b011100111011101110: begin rgb_reg = 3'b111; end
            18'b011100111011110001: begin rgb_reg = 3'b111; end
            18'b011100111011110010: begin rgb_reg = 3'b111; end
            18'b011100111011110101: begin rgb_reg = 3'b111; end
            18'b011100111011110110: begin rgb_reg = 3'b111; end
            18'b011100111011111011: begin rgb_reg = 3'b111; end
            18'b011100111011111100: begin rgb_reg = 3'b111; end
            18'b011100111011111101: begin rgb_reg = 3'b111; end
            18'b011100111011111110: begin rgb_reg = 3'b111; end
            18'b011100111011111111: begin rgb_reg = 3'b111; end
            18'b011100111100000000: begin rgb_reg = 3'b111; end
            18'b011100111100000111: begin rgb_reg = 3'b111; end
            18'b011100111100001000: begin rgb_reg = 3'b111; end
            18'b011100111100001101: begin rgb_reg = 3'b111; end
            18'b011100111100001110: begin rgb_reg = 3'b111; end
            18'b011100111100010001: begin rgb_reg = 3'b111; end
            18'b011100111100010010: begin rgb_reg = 3'b111; end
            18'b011100111100010011: begin rgb_reg = 3'b111; end
            18'b011100111100010100: begin rgb_reg = 3'b111; end
            18'b011100111100011011: begin rgb_reg = 3'b111; end
            18'b011100111100011100: begin rgb_reg = 3'b111; end
            18'b011100111100011101: begin rgb_reg = 3'b111; end
            18'b011100111100011110: begin rgb_reg = 3'b111; end
            18'b011100111100011111: begin rgb_reg = 3'b111; end
            18'b011100111100100000: begin rgb_reg = 3'b111; end
            18'b011100111100100111: begin rgb_reg = 3'b111; end
            18'b011100111100101000: begin rgb_reg = 3'b111; end
            18'b011100111100101001: begin rgb_reg = 3'b111; end
            18'b011100111100101010: begin rgb_reg = 3'b111; end
            18'b011100111100101011: begin rgb_reg = 3'b111; end
            18'b011100111100101100: begin rgb_reg = 3'b111; end
            18'b011100111100101101: begin rgb_reg = 3'b111; end
            18'b011100111100101110: begin rgb_reg = 3'b111; end
            18'b011100111100110011: begin rgb_reg = 3'b111; end
            18'b011100111100110100: begin rgb_reg = 3'b111; end
            18'b011100111100110101: begin rgb_reg = 3'b111; end
            18'b011100111100110110: begin rgb_reg = 3'b111; end
            18'b011100111100110111: begin rgb_reg = 3'b111; end
            18'b011100111100111000: begin rgb_reg = 3'b111; end
            18'b011100111100111111: begin rgb_reg = 3'b111; end
            18'b011100111101000000: begin rgb_reg = 3'b111; end
            18'b011100111101000111: begin rgb_reg = 3'b111; end
            18'b011100111101001000: begin rgb_reg = 3'b111; end
            18'b011100111101001001: begin rgb_reg = 3'b111; end
            18'b011100111101001010: begin rgb_reg = 3'b111; end
            18'b011100111101001011: begin rgb_reg = 3'b111; end
            18'b011100111101001100: begin rgb_reg = 3'b111; end
            18'b011101000010110001: begin rgb_reg = 3'b111; end
            18'b011101000010110010: begin rgb_reg = 3'b111; end
            18'b011101000010111001: begin rgb_reg = 3'b111; end
            18'b011101000010111010: begin rgb_reg = 3'b111; end
            18'b011101000010111101: begin rgb_reg = 3'b111; end
            18'b011101000010111110: begin rgb_reg = 3'b111; end
            18'b011101000011000101: begin rgb_reg = 3'b111; end
            18'b011101000011000110: begin rgb_reg = 3'b111; end
            18'b011101000011010001: begin rgb_reg = 3'b111; end
            18'b011101000011010010: begin rgb_reg = 3'b111; end
            18'b011101000011010101: begin rgb_reg = 3'b111; end
            18'b011101000011010110: begin rgb_reg = 3'b111; end
            18'b011101000011011101: begin rgb_reg = 3'b111; end
            18'b011101000011011110: begin rgb_reg = 3'b111; end
            18'b011101000011101101: begin rgb_reg = 3'b111; end
            18'b011101000011101110: begin rgb_reg = 3'b111; end
            18'b011101000011110101: begin rgb_reg = 3'b111; end
            18'b011101000011110110: begin rgb_reg = 3'b111; end
            18'b011101000011111001: begin rgb_reg = 3'b111; end
            18'b011101000011111010: begin rgb_reg = 3'b111; end
            18'b011101000100000001: begin rgb_reg = 3'b111; end
            18'b011101000100000010: begin rgb_reg = 3'b111; end
            18'b011101000100000111: begin rgb_reg = 3'b111; end
            18'b011101000100001000: begin rgb_reg = 3'b111; end
            18'b011101000100001101: begin rgb_reg = 3'b111; end
            18'b011101000100001110: begin rgb_reg = 3'b111; end
            18'b011101000100001111: begin rgb_reg = 3'b111; end
            18'b011101000100010000: begin rgb_reg = 3'b111; end
            18'b011101000100010101: begin rgb_reg = 3'b111; end
            18'b011101000100010110: begin rgb_reg = 3'b111; end
            18'b011101000100100001: begin rgb_reg = 3'b111; end
            18'b011101000100100010: begin rgb_reg = 3'b111; end
            18'b011101000100100101: begin rgb_reg = 3'b111; end
            18'b011101000100100110: begin rgb_reg = 3'b111; end
            18'b011101000100111001: begin rgb_reg = 3'b111; end
            18'b011101000100111010: begin rgb_reg = 3'b111; end
            18'b011101000100111111: begin rgb_reg = 3'b111; end
            18'b011101000101000000: begin rgb_reg = 3'b111; end
            18'b011101000101000101: begin rgb_reg = 3'b111; end
            18'b011101000101000110: begin rgb_reg = 3'b111; end
            18'b011101000101001101: begin rgb_reg = 3'b111; end
            18'b011101000101001110: begin rgb_reg = 3'b111; end
            18'b011101001010110001: begin rgb_reg = 3'b111; end
            18'b011101001010110010: begin rgb_reg = 3'b111; end
            18'b011101001010111001: begin rgb_reg = 3'b111; end
            18'b011101001010111010: begin rgb_reg = 3'b111; end
            18'b011101001010111101: begin rgb_reg = 3'b111; end
            18'b011101001010111110: begin rgb_reg = 3'b111; end
            18'b011101001011000101: begin rgb_reg = 3'b111; end
            18'b011101001011000110: begin rgb_reg = 3'b111; end
            18'b011101001011010001: begin rgb_reg = 3'b111; end
            18'b011101001011010010: begin rgb_reg = 3'b111; end
            18'b011101001011010101: begin rgb_reg = 3'b111; end
            18'b011101001011010110: begin rgb_reg = 3'b111; end
            18'b011101001011011101: begin rgb_reg = 3'b111; end
            18'b011101001011011110: begin rgb_reg = 3'b111; end
            18'b011101001011101101: begin rgb_reg = 3'b111; end
            18'b011101001011101110: begin rgb_reg = 3'b111; end
            18'b011101001011110101: begin rgb_reg = 3'b111; end
            18'b011101001011110110: begin rgb_reg = 3'b111; end
            18'b011101001011111001: begin rgb_reg = 3'b111; end
            18'b011101001011111010: begin rgb_reg = 3'b111; end
            18'b011101001100000001: begin rgb_reg = 3'b111; end
            18'b011101001100000010: begin rgb_reg = 3'b111; end
            18'b011101001100000111: begin rgb_reg = 3'b111; end
            18'b011101001100001000: begin rgb_reg = 3'b111; end
            18'b011101001100001101: begin rgb_reg = 3'b111; end
            18'b011101001100001110: begin rgb_reg = 3'b111; end
            18'b011101001100001111: begin rgb_reg = 3'b111; end
            18'b011101001100010000: begin rgb_reg = 3'b111; end
            18'b011101001100010101: begin rgb_reg = 3'b111; end
            18'b011101001100010110: begin rgb_reg = 3'b111; end
            18'b011101001100100001: begin rgb_reg = 3'b111; end
            18'b011101001100100010: begin rgb_reg = 3'b111; end
            18'b011101001100100101: begin rgb_reg = 3'b111; end
            18'b011101001100100110: begin rgb_reg = 3'b111; end
            18'b011101001100111001: begin rgb_reg = 3'b111; end
            18'b011101001100111010: begin rgb_reg = 3'b111; end
            18'b011101001100111111: begin rgb_reg = 3'b111; end
            18'b011101001101000000: begin rgb_reg = 3'b111; end
            18'b011101001101000101: begin rgb_reg = 3'b111; end
            18'b011101001101000110: begin rgb_reg = 3'b111; end
            18'b011101001101001101: begin rgb_reg = 3'b111; end
            18'b011101001101001110: begin rgb_reg = 3'b111; end
            18'b011101010010110001: begin rgb_reg = 3'b111; end
            18'b011101010010110010: begin rgb_reg = 3'b111; end
            18'b011101010010111001: begin rgb_reg = 3'b111; end
            18'b011101010010111010: begin rgb_reg = 3'b111; end
            18'b011101010010111101: begin rgb_reg = 3'b111; end
            18'b011101010010111110: begin rgb_reg = 3'b111; end
            18'b011101010011000101: begin rgb_reg = 3'b111; end
            18'b011101010011000110: begin rgb_reg = 3'b111; end
            18'b011101010011001011: begin rgb_reg = 3'b111; end
            18'b011101010011001100: begin rgb_reg = 3'b111; end
            18'b011101010011001101: begin rgb_reg = 3'b111; end
            18'b011101010011001110: begin rgb_reg = 3'b111; end
            18'b011101010011001111: begin rgb_reg = 3'b111; end
            18'b011101010011010000: begin rgb_reg = 3'b111; end
            18'b011101010011010001: begin rgb_reg = 3'b111; end
            18'b011101010011010010: begin rgb_reg = 3'b111; end
            18'b011101010011010101: begin rgb_reg = 3'b111; end
            18'b011101010011010110: begin rgb_reg = 3'b111; end
            18'b011101010011011101: begin rgb_reg = 3'b111; end
            18'b011101010011011110: begin rgb_reg = 3'b111; end
            18'b011101010011101101: begin rgb_reg = 3'b111; end
            18'b011101010011101110: begin rgb_reg = 3'b111; end
            18'b011101010011110101: begin rgb_reg = 3'b111; end
            18'b011101010011110110: begin rgb_reg = 3'b111; end
            18'b011101010011111001: begin rgb_reg = 3'b111; end
            18'b011101010011111010: begin rgb_reg = 3'b111; end
            18'b011101010011111011: begin rgb_reg = 3'b111; end
            18'b011101010011111100: begin rgb_reg = 3'b111; end
            18'b011101010011111101: begin rgb_reg = 3'b111; end
            18'b011101010011111110: begin rgb_reg = 3'b111; end
            18'b011101010011111111: begin rgb_reg = 3'b111; end
            18'b011101010100000000: begin rgb_reg = 3'b111; end
            18'b011101010100000001: begin rgb_reg = 3'b111; end
            18'b011101010100000010: begin rgb_reg = 3'b111; end
            18'b011101010100000111: begin rgb_reg = 3'b111; end
            18'b011101010100001000: begin rgb_reg = 3'b111; end
            18'b011101010100001101: begin rgb_reg = 3'b111; end
            18'b011101010100001110: begin rgb_reg = 3'b111; end
            18'b011101010100010101: begin rgb_reg = 3'b111; end
            18'b011101010100010110: begin rgb_reg = 3'b111; end
            18'b011101010100011011: begin rgb_reg = 3'b111; end
            18'b011101010100011100: begin rgb_reg = 3'b111; end
            18'b011101010100011101: begin rgb_reg = 3'b111; end
            18'b011101010100011110: begin rgb_reg = 3'b111; end
            18'b011101010100011111: begin rgb_reg = 3'b111; end
            18'b011101010100100000: begin rgb_reg = 3'b111; end
            18'b011101010100100001: begin rgb_reg = 3'b111; end
            18'b011101010100100010: begin rgb_reg = 3'b111; end
            18'b011101010100100111: begin rgb_reg = 3'b111; end
            18'b011101010100101000: begin rgb_reg = 3'b111; end
            18'b011101010100101001: begin rgb_reg = 3'b111; end
            18'b011101010100101010: begin rgb_reg = 3'b111; end
            18'b011101010100101011: begin rgb_reg = 3'b111; end
            18'b011101010100101100: begin rgb_reg = 3'b111; end
            18'b011101010100110011: begin rgb_reg = 3'b111; end
            18'b011101010100110100: begin rgb_reg = 3'b111; end
            18'b011101010100110101: begin rgb_reg = 3'b111; end
            18'b011101010100110110: begin rgb_reg = 3'b111; end
            18'b011101010100110111: begin rgb_reg = 3'b111; end
            18'b011101010100111000: begin rgb_reg = 3'b111; end
            18'b011101010100111001: begin rgb_reg = 3'b111; end
            18'b011101010100111010: begin rgb_reg = 3'b111; end
            18'b011101010100111111: begin rgb_reg = 3'b111; end
            18'b011101010101000000: begin rgb_reg = 3'b111; end
            18'b011101010101000101: begin rgb_reg = 3'b111; end
            18'b011101010101000110: begin rgb_reg = 3'b111; end
            18'b011101010101000111: begin rgb_reg = 3'b111; end
            18'b011101010101001000: begin rgb_reg = 3'b111; end
            18'b011101010101001001: begin rgb_reg = 3'b111; end
            18'b011101010101001010: begin rgb_reg = 3'b111; end
            18'b011101010101001011: begin rgb_reg = 3'b111; end
            18'b011101010101001100: begin rgb_reg = 3'b111; end
            18'b011101010101001101: begin rgb_reg = 3'b111; end
            18'b011101010101001110: begin rgb_reg = 3'b111; end
            18'b011101011010110001: begin rgb_reg = 3'b111; end
            18'b011101011010110010: begin rgb_reg = 3'b111; end
            18'b011101011010111001: begin rgb_reg = 3'b111; end
            18'b011101011010111010: begin rgb_reg = 3'b111; end
            18'b011101011010111101: begin rgb_reg = 3'b111; end
            18'b011101011010111110: begin rgb_reg = 3'b111; end
            18'b011101011011000101: begin rgb_reg = 3'b111; end
            18'b011101011011000110: begin rgb_reg = 3'b111; end
            18'b011101011011001011: begin rgb_reg = 3'b111; end
            18'b011101011011001100: begin rgb_reg = 3'b111; end
            18'b011101011011001101: begin rgb_reg = 3'b111; end
            18'b011101011011001110: begin rgb_reg = 3'b111; end
            18'b011101011011001111: begin rgb_reg = 3'b111; end
            18'b011101011011010000: begin rgb_reg = 3'b111; end
            18'b011101011011010001: begin rgb_reg = 3'b111; end
            18'b011101011011010010: begin rgb_reg = 3'b111; end
            18'b011101011011010101: begin rgb_reg = 3'b111; end
            18'b011101011011010110: begin rgb_reg = 3'b111; end
            18'b011101011011011101: begin rgb_reg = 3'b111; end
            18'b011101011011011110: begin rgb_reg = 3'b111; end
            18'b011101011011101101: begin rgb_reg = 3'b111; end
            18'b011101011011101110: begin rgb_reg = 3'b111; end
            18'b011101011011110101: begin rgb_reg = 3'b111; end
            18'b011101011011110110: begin rgb_reg = 3'b111; end
            18'b011101011011111001: begin rgb_reg = 3'b111; end
            18'b011101011011111010: begin rgb_reg = 3'b111; end
            18'b011101011011111011: begin rgb_reg = 3'b111; end
            18'b011101011011111100: begin rgb_reg = 3'b111; end
            18'b011101011011111101: begin rgb_reg = 3'b111; end
            18'b011101011011111110: begin rgb_reg = 3'b111; end
            18'b011101011011111111: begin rgb_reg = 3'b111; end
            18'b011101011100000000: begin rgb_reg = 3'b111; end
            18'b011101011100000001: begin rgb_reg = 3'b111; end
            18'b011101011100000010: begin rgb_reg = 3'b111; end
            18'b011101011100000111: begin rgb_reg = 3'b111; end
            18'b011101011100001000: begin rgb_reg = 3'b111; end
            18'b011101011100001101: begin rgb_reg = 3'b111; end
            18'b011101011100001110: begin rgb_reg = 3'b111; end
            18'b011101011100010101: begin rgb_reg = 3'b111; end
            18'b011101011100010110: begin rgb_reg = 3'b111; end
            18'b011101011100011011: begin rgb_reg = 3'b111; end
            18'b011101011100011100: begin rgb_reg = 3'b111; end
            18'b011101011100011101: begin rgb_reg = 3'b111; end
            18'b011101011100011110: begin rgb_reg = 3'b111; end
            18'b011101011100011111: begin rgb_reg = 3'b111; end
            18'b011101011100100000: begin rgb_reg = 3'b111; end
            18'b011101011100100001: begin rgb_reg = 3'b111; end
            18'b011101011100100010: begin rgb_reg = 3'b111; end
            18'b011101011100100111: begin rgb_reg = 3'b111; end
            18'b011101011100101000: begin rgb_reg = 3'b111; end
            18'b011101011100101001: begin rgb_reg = 3'b111; end
            18'b011101011100101010: begin rgb_reg = 3'b111; end
            18'b011101011100101011: begin rgb_reg = 3'b111; end
            18'b011101011100101100: begin rgb_reg = 3'b111; end
            18'b011101011100110011: begin rgb_reg = 3'b111; end
            18'b011101011100110100: begin rgb_reg = 3'b111; end
            18'b011101011100110101: begin rgb_reg = 3'b111; end
            18'b011101011100110110: begin rgb_reg = 3'b111; end
            18'b011101011100110111: begin rgb_reg = 3'b111; end
            18'b011101011100111000: begin rgb_reg = 3'b111; end
            18'b011101011100111001: begin rgb_reg = 3'b111; end
            18'b011101011100111010: begin rgb_reg = 3'b111; end
            18'b011101011100111111: begin rgb_reg = 3'b111; end
            18'b011101011101000000: begin rgb_reg = 3'b111; end
            18'b011101011101000101: begin rgb_reg = 3'b111; end
            18'b011101011101000110: begin rgb_reg = 3'b111; end
            18'b011101011101000111: begin rgb_reg = 3'b111; end
            18'b011101011101001000: begin rgb_reg = 3'b111; end
            18'b011101011101001001: begin rgb_reg = 3'b111; end
            18'b011101011101001010: begin rgb_reg = 3'b111; end
            18'b011101011101001011: begin rgb_reg = 3'b111; end
            18'b011101011101001100: begin rgb_reg = 3'b111; end
            18'b011101011101001101: begin rgb_reg = 3'b111; end
            18'b011101011101001110: begin rgb_reg = 3'b111; end
            18'b011101100010110001: begin rgb_reg = 3'b111; end
            18'b011101100010110010: begin rgb_reg = 3'b111; end
            18'b011101100010111001: begin rgb_reg = 3'b111; end
            18'b011101100010111010: begin rgb_reg = 3'b111; end
            18'b011101100010111101: begin rgb_reg = 3'b111; end
            18'b011101100010111110: begin rgb_reg = 3'b111; end
            18'b011101100011000101: begin rgb_reg = 3'b111; end
            18'b011101100011000110: begin rgb_reg = 3'b111; end
            18'b011101100011001001: begin rgb_reg = 3'b111; end
            18'b011101100011001010: begin rgb_reg = 3'b111; end
            18'b011101100011010001: begin rgb_reg = 3'b111; end
            18'b011101100011010010: begin rgb_reg = 3'b111; end
            18'b011101100011010101: begin rgb_reg = 3'b111; end
            18'b011101100011010110: begin rgb_reg = 3'b111; end
            18'b011101100011011101: begin rgb_reg = 3'b111; end
            18'b011101100011011110: begin rgb_reg = 3'b111; end
            18'b011101100011101101: begin rgb_reg = 3'b111; end
            18'b011101100011101110: begin rgb_reg = 3'b111; end
            18'b011101100011110101: begin rgb_reg = 3'b111; end
            18'b011101100011110110: begin rgb_reg = 3'b111; end
            18'b011101100011111001: begin rgb_reg = 3'b111; end
            18'b011101100011111010: begin rgb_reg = 3'b111; end
            18'b011101100100000111: begin rgb_reg = 3'b111; end
            18'b011101100100001000: begin rgb_reg = 3'b111; end
            18'b011101100100001101: begin rgb_reg = 3'b111; end
            18'b011101100100001110: begin rgb_reg = 3'b111; end
            18'b011101100100010101: begin rgb_reg = 3'b111; end
            18'b011101100100010110: begin rgb_reg = 3'b111; end
            18'b011101100100011001: begin rgb_reg = 3'b111; end
            18'b011101100100011010: begin rgb_reg = 3'b111; end
            18'b011101100100100001: begin rgb_reg = 3'b111; end
            18'b011101100100100010: begin rgb_reg = 3'b111; end
            18'b011101100100101101: begin rgb_reg = 3'b111; end
            18'b011101100100101110: begin rgb_reg = 3'b111; end
            18'b011101100100110001: begin rgb_reg = 3'b111; end
            18'b011101100100110010: begin rgb_reg = 3'b111; end
            18'b011101100100111001: begin rgb_reg = 3'b111; end
            18'b011101100100111010: begin rgb_reg = 3'b111; end
            18'b011101100100111111: begin rgb_reg = 3'b111; end
            18'b011101100101000000: begin rgb_reg = 3'b111; end
            18'b011101100101000101: begin rgb_reg = 3'b111; end
            18'b011101100101000110: begin rgb_reg = 3'b111; end
            18'b011101101010110001: begin rgb_reg = 3'b111; end
            18'b011101101010110010: begin rgb_reg = 3'b111; end
            18'b011101101010111001: begin rgb_reg = 3'b111; end
            18'b011101101010111010: begin rgb_reg = 3'b111; end
            18'b011101101010111101: begin rgb_reg = 3'b111; end
            18'b011101101010111110: begin rgb_reg = 3'b111; end
            18'b011101101011000101: begin rgb_reg = 3'b111; end
            18'b011101101011000110: begin rgb_reg = 3'b111; end
            18'b011101101011001001: begin rgb_reg = 3'b111; end
            18'b011101101011001010: begin rgb_reg = 3'b111; end
            18'b011101101011010001: begin rgb_reg = 3'b111; end
            18'b011101101011010010: begin rgb_reg = 3'b111; end
            18'b011101101011010101: begin rgb_reg = 3'b111; end
            18'b011101101011010110: begin rgb_reg = 3'b111; end
            18'b011101101011011101: begin rgb_reg = 3'b111; end
            18'b011101101011011110: begin rgb_reg = 3'b111; end
            18'b011101101011101101: begin rgb_reg = 3'b111; end
            18'b011101101011101110: begin rgb_reg = 3'b111; end
            18'b011101101011110101: begin rgb_reg = 3'b111; end
            18'b011101101011110110: begin rgb_reg = 3'b111; end
            18'b011101101011111001: begin rgb_reg = 3'b111; end
            18'b011101101011111010: begin rgb_reg = 3'b111; end
            18'b011101101100000111: begin rgb_reg = 3'b111; end
            18'b011101101100001000: begin rgb_reg = 3'b111; end
            18'b011101101100001101: begin rgb_reg = 3'b111; end
            18'b011101101100001110: begin rgb_reg = 3'b111; end
            18'b011101101100010101: begin rgb_reg = 3'b111; end
            18'b011101101100010110: begin rgb_reg = 3'b111; end
            18'b011101101100011001: begin rgb_reg = 3'b111; end
            18'b011101101100011010: begin rgb_reg = 3'b111; end
            18'b011101101100100001: begin rgb_reg = 3'b111; end
            18'b011101101100100010: begin rgb_reg = 3'b111; end
            18'b011101101100101101: begin rgb_reg = 3'b111; end
            18'b011101101100101110: begin rgb_reg = 3'b111; end
            18'b011101101100110001: begin rgb_reg = 3'b111; end
            18'b011101101100110010: begin rgb_reg = 3'b111; end
            18'b011101101100111001: begin rgb_reg = 3'b111; end
            18'b011101101100111010: begin rgb_reg = 3'b111; end
            18'b011101101100111111: begin rgb_reg = 3'b111; end
            18'b011101101101000000: begin rgb_reg = 3'b111; end
            18'b011101101101000101: begin rgb_reg = 3'b111; end
            18'b011101101101000110: begin rgb_reg = 3'b111; end
            18'b011101110010110001: begin rgb_reg = 3'b111; end
            18'b011101110010110010: begin rgb_reg = 3'b111; end
            18'b011101110010111001: begin rgb_reg = 3'b111; end
            18'b011101110010111010: begin rgb_reg = 3'b111; end
            18'b011101110010111101: begin rgb_reg = 3'b111; end
            18'b011101110010111110: begin rgb_reg = 3'b111; end
            18'b011101110011000101: begin rgb_reg = 3'b111; end
            18'b011101110011000110: begin rgb_reg = 3'b111; end
            18'b011101110011001011: begin rgb_reg = 3'b111; end
            18'b011101110011001100: begin rgb_reg = 3'b111; end
            18'b011101110011001101: begin rgb_reg = 3'b111; end
            18'b011101110011001110: begin rgb_reg = 3'b111; end
            18'b011101110011001111: begin rgb_reg = 3'b111; end
            18'b011101110011010000: begin rgb_reg = 3'b111; end
            18'b011101110011010001: begin rgb_reg = 3'b111; end
            18'b011101110011010010: begin rgb_reg = 3'b111; end
            18'b011101110011010101: begin rgb_reg = 3'b111; end
            18'b011101110011010110: begin rgb_reg = 3'b111; end
            18'b011101110011011101: begin rgb_reg = 3'b111; end
            18'b011101110011011110: begin rgb_reg = 3'b111; end
            18'b011101110011101101: begin rgb_reg = 3'b111; end
            18'b011101110011101110: begin rgb_reg = 3'b111; end
            18'b011101110011110101: begin rgb_reg = 3'b111; end
            18'b011101110011110110: begin rgb_reg = 3'b111; end
            18'b011101110011111011: begin rgb_reg = 3'b111; end
            18'b011101110011111100: begin rgb_reg = 3'b111; end
            18'b011101110011111101: begin rgb_reg = 3'b111; end
            18'b011101110011111110: begin rgb_reg = 3'b111; end
            18'b011101110011111111: begin rgb_reg = 3'b111; end
            18'b011101110100000000: begin rgb_reg = 3'b111; end
            18'b011101110100000001: begin rgb_reg = 3'b111; end
            18'b011101110100000010: begin rgb_reg = 3'b111; end
            18'b011101110100001001: begin rgb_reg = 3'b111; end
            18'b011101110100001010: begin rgb_reg = 3'b111; end
            18'b011101110100001101: begin rgb_reg = 3'b111; end
            18'b011101110100001110: begin rgb_reg = 3'b111; end
            18'b011101110100010101: begin rgb_reg = 3'b111; end
            18'b011101110100010110: begin rgb_reg = 3'b111; end
            18'b011101110100011011: begin rgb_reg = 3'b111; end
            18'b011101110100011100: begin rgb_reg = 3'b111; end
            18'b011101110100011101: begin rgb_reg = 3'b111; end
            18'b011101110100011110: begin rgb_reg = 3'b111; end
            18'b011101110100011111: begin rgb_reg = 3'b111; end
            18'b011101110100100000: begin rgb_reg = 3'b111; end
            18'b011101110100100001: begin rgb_reg = 3'b111; end
            18'b011101110100100010: begin rgb_reg = 3'b111; end
            18'b011101110100100101: begin rgb_reg = 3'b111; end
            18'b011101110100100110: begin rgb_reg = 3'b111; end
            18'b011101110100100111: begin rgb_reg = 3'b111; end
            18'b011101110100101000: begin rgb_reg = 3'b111; end
            18'b011101110100101001: begin rgb_reg = 3'b111; end
            18'b011101110100101010: begin rgb_reg = 3'b111; end
            18'b011101110100101011: begin rgb_reg = 3'b111; end
            18'b011101110100101100: begin rgb_reg = 3'b111; end
            18'b011101110100110011: begin rgb_reg = 3'b111; end
            18'b011101110100110100: begin rgb_reg = 3'b111; end
            18'b011101110100110101: begin rgb_reg = 3'b111; end
            18'b011101110100110110: begin rgb_reg = 3'b111; end
            18'b011101110100110111: begin rgb_reg = 3'b111; end
            18'b011101110100111000: begin rgb_reg = 3'b111; end
            18'b011101110100111001: begin rgb_reg = 3'b111; end
            18'b011101110100111010: begin rgb_reg = 3'b111; end
            18'b011101110101000001: begin rgb_reg = 3'b111; end
            18'b011101110101000010: begin rgb_reg = 3'b111; end
            18'b011101110101000111: begin rgb_reg = 3'b111; end
            18'b011101110101001000: begin rgb_reg = 3'b111; end
            18'b011101110101001001: begin rgb_reg = 3'b111; end
            18'b011101110101001010: begin rgb_reg = 3'b111; end
            18'b011101110101001011: begin rgb_reg = 3'b111; end
            18'b011101110101001100: begin rgb_reg = 3'b111; end
            18'b011101110101001101: begin rgb_reg = 3'b111; end
            18'b011101110101001110: begin rgb_reg = 3'b111; end
            18'b011101111010110001: begin rgb_reg = 3'b111; end
            18'b011101111010110010: begin rgb_reg = 3'b111; end
            18'b011101111010111001: begin rgb_reg = 3'b111; end
            18'b011101111010111010: begin rgb_reg = 3'b111; end
            18'b011101111010111101: begin rgb_reg = 3'b111; end
            18'b011101111010111110: begin rgb_reg = 3'b111; end
            18'b011101111011000101: begin rgb_reg = 3'b111; end
            18'b011101111011000110: begin rgb_reg = 3'b111; end
            18'b011101111011001011: begin rgb_reg = 3'b111; end
            18'b011101111011001100: begin rgb_reg = 3'b111; end
            18'b011101111011001101: begin rgb_reg = 3'b111; end
            18'b011101111011001110: begin rgb_reg = 3'b111; end
            18'b011101111011001111: begin rgb_reg = 3'b111; end
            18'b011101111011010000: begin rgb_reg = 3'b111; end
            18'b011101111011010001: begin rgb_reg = 3'b111; end
            18'b011101111011010010: begin rgb_reg = 3'b111; end
            18'b011101111011010101: begin rgb_reg = 3'b111; end
            18'b011101111011010110: begin rgb_reg = 3'b111; end
            18'b011101111011011101: begin rgb_reg = 3'b111; end
            18'b011101111011011110: begin rgb_reg = 3'b111; end
            18'b011101111011101101: begin rgb_reg = 3'b111; end
            18'b011101111011101110: begin rgb_reg = 3'b111; end
            18'b011101111011110101: begin rgb_reg = 3'b111; end
            18'b011101111011110110: begin rgb_reg = 3'b111; end
            18'b011101111011111011: begin rgb_reg = 3'b111; end
            18'b011101111011111100: begin rgb_reg = 3'b111; end
            18'b011101111011111101: begin rgb_reg = 3'b111; end
            18'b011101111011111110: begin rgb_reg = 3'b111; end
            18'b011101111011111111: begin rgb_reg = 3'b111; end
            18'b011101111100000000: begin rgb_reg = 3'b111; end
            18'b011101111100000001: begin rgb_reg = 3'b111; end
            18'b011101111100000010: begin rgb_reg = 3'b111; end
            18'b011101111100001001: begin rgb_reg = 3'b111; end
            18'b011101111100001010: begin rgb_reg = 3'b111; end
            18'b011101111100001101: begin rgb_reg = 3'b111; end
            18'b011101111100001110: begin rgb_reg = 3'b111; end
            18'b011101111100010101: begin rgb_reg = 3'b111; end
            18'b011101111100010110: begin rgb_reg = 3'b111; end
            18'b011101111100011011: begin rgb_reg = 3'b111; end
            18'b011101111100011100: begin rgb_reg = 3'b111; end
            18'b011101111100011101: begin rgb_reg = 3'b111; end
            18'b011101111100011110: begin rgb_reg = 3'b111; end
            18'b011101111100011111: begin rgb_reg = 3'b111; end
            18'b011101111100100000: begin rgb_reg = 3'b111; end
            18'b011101111100100001: begin rgb_reg = 3'b111; end
            18'b011101111100100010: begin rgb_reg = 3'b111; end
            18'b011101111100100101: begin rgb_reg = 3'b111; end
            18'b011101111100100110: begin rgb_reg = 3'b111; end
            18'b011101111100100111: begin rgb_reg = 3'b111; end
            18'b011101111100101000: begin rgb_reg = 3'b111; end
            18'b011101111100101001: begin rgb_reg = 3'b111; end
            18'b011101111100101010: begin rgb_reg = 3'b111; end
            18'b011101111100101011: begin rgb_reg = 3'b111; end
            18'b011101111100101100: begin rgb_reg = 3'b111; end
            18'b011101111100110011: begin rgb_reg = 3'b111; end
            18'b011101111100110100: begin rgb_reg = 3'b111; end
            18'b011101111100110101: begin rgb_reg = 3'b111; end
            18'b011101111100110110: begin rgb_reg = 3'b111; end
            18'b011101111100110111: begin rgb_reg = 3'b111; end
            18'b011101111100111000: begin rgb_reg = 3'b111; end
            18'b011101111100111001: begin rgb_reg = 3'b111; end
            18'b011101111100111010: begin rgb_reg = 3'b111; end
            18'b011101111101000001: begin rgb_reg = 3'b111; end
            18'b011101111101000010: begin rgb_reg = 3'b111; end
            18'b011101111101000111: begin rgb_reg = 3'b111; end
            18'b011101111101001000: begin rgb_reg = 3'b111; end
            18'b011101111101001001: begin rgb_reg = 3'b111; end
            18'b011101111101001010: begin rgb_reg = 3'b111; end
            18'b011101111101001011: begin rgb_reg = 3'b111; end
            18'b011101111101001100: begin rgb_reg = 3'b111; end
            18'b011101111101001101: begin rgb_reg = 3'b111; end
            18'b011101111101001110: begin rgb_reg = 3'b111; end
            18'b100000101011000010: begin rgb_reg = 3'b111; end
            18'b100000101011000011: begin rgb_reg = 3'b111; end
            18'b100000101011000100: begin rgb_reg = 3'b111; end
            18'b100000101011000101: begin rgb_reg = 3'b111; end
            18'b100000101011000110: begin rgb_reg = 3'b111; end
            18'b100000101011001101: begin rgb_reg = 3'b111; end
            18'b100000101011001110: begin rgb_reg = 3'b111; end
            18'b100000101011001111: begin rgb_reg = 3'b111; end
            18'b100000101011010000: begin rgb_reg = 3'b111; end
            18'b100000101011010001: begin rgb_reg = 3'b111; end
            18'b100000101011010010: begin rgb_reg = 3'b111; end
            18'b100000101011010011: begin rgb_reg = 3'b111; end
            18'b100000101011011011: begin rgb_reg = 3'b111; end
            18'b100000101011011100: begin rgb_reg = 3'b111; end
            18'b100000101011011101: begin rgb_reg = 3'b111; end
            18'b100000101011011110: begin rgb_reg = 3'b111; end
            18'b100000101011011111: begin rgb_reg = 3'b111; end
            18'b100000101011100000: begin rgb_reg = 3'b111; end
            18'b100000101011100001: begin rgb_reg = 3'b111; end
            18'b100000101011101000: begin rgb_reg = 3'b111; end
            18'b100000101011101001: begin rgb_reg = 3'b111; end
            18'b100000101011101010: begin rgb_reg = 3'b111; end
            18'b100000101011101011: begin rgb_reg = 3'b111; end
            18'b100000101011101100: begin rgb_reg = 3'b111; end
            18'b100000101011101101: begin rgb_reg = 3'b111; end
            18'b100000101011101110: begin rgb_reg = 3'b111; end
            18'b100000101011110110: begin rgb_reg = 3'b111; end
            18'b100000101011110111: begin rgb_reg = 3'b111; end
            18'b100000101011111000: begin rgb_reg = 3'b111; end
            18'b100000101011111001: begin rgb_reg = 3'b111; end
            18'b100000101011111010: begin rgb_reg = 3'b111; end
            18'b100000101011111011: begin rgb_reg = 3'b111; end
            18'b100000101011111100: begin rgb_reg = 3'b111; end
            18'b100000101100000011: begin rgb_reg = 3'b111; end
            18'b100000101100000100: begin rgb_reg = 3'b111; end
            18'b100000101100000101: begin rgb_reg = 3'b111; end
            18'b100000101100000110: begin rgb_reg = 3'b111; end
            18'b100000101100000111: begin rgb_reg = 3'b111; end
            18'b100000101100001000: begin rgb_reg = 3'b111; end
            18'b100000101100001001: begin rgb_reg = 3'b111; end
            18'b100000101100010011: begin rgb_reg = 3'b111; end
            18'b100000101100010100: begin rgb_reg = 3'b111; end
            18'b100000101100010101: begin rgb_reg = 3'b111; end
            18'b100000101100010110: begin rgb_reg = 3'b111; end
            18'b100000101100010111: begin rgb_reg = 3'b111; end
            18'b100000101100100001: begin rgb_reg = 3'b111; end
            18'b100000101100100010: begin rgb_reg = 3'b111; end
            18'b100000101100101100: begin rgb_reg = 3'b111; end
            18'b100000101100101101: begin rgb_reg = 3'b111; end
            18'b100000101100101110: begin rgb_reg = 3'b111; end
            18'b100000101100101111: begin rgb_reg = 3'b111; end
            18'b100000101100110000: begin rgb_reg = 3'b111; end
            18'b100000101100110001: begin rgb_reg = 3'b111; end
            18'b100000101100110010: begin rgb_reg = 3'b111; end
            18'b100000101100111100: begin rgb_reg = 3'b111; end
            18'b100000101100111101: begin rgb_reg = 3'b111; end
            18'b100000110011000010: begin rgb_reg = 3'b111; end
            18'b100000110011000011: begin rgb_reg = 3'b111; end
            18'b100000110011000100: begin rgb_reg = 3'b111; end
            18'b100000110011000101: begin rgb_reg = 3'b111; end
            18'b100000110011000110: begin rgb_reg = 3'b111; end
            18'b100000110011001101: begin rgb_reg = 3'b111; end
            18'b100000110011001110: begin rgb_reg = 3'b111; end
            18'b100000110011001111: begin rgb_reg = 3'b111; end
            18'b100000110011010000: begin rgb_reg = 3'b111; end
            18'b100000110011010001: begin rgb_reg = 3'b111; end
            18'b100000110011010010: begin rgb_reg = 3'b111; end
            18'b100000110011010011: begin rgb_reg = 3'b111; end
            18'b100000110011011011: begin rgb_reg = 3'b111; end
            18'b100000110011011100: begin rgb_reg = 3'b111; end
            18'b100000110011011101: begin rgb_reg = 3'b111; end
            18'b100000110011011110: begin rgb_reg = 3'b111; end
            18'b100000110011011111: begin rgb_reg = 3'b111; end
            18'b100000110011100000: begin rgb_reg = 3'b111; end
            18'b100000110011100001: begin rgb_reg = 3'b111; end
            18'b100000110011101000: begin rgb_reg = 3'b111; end
            18'b100000110011101001: begin rgb_reg = 3'b111; end
            18'b100000110011101010: begin rgb_reg = 3'b111; end
            18'b100000110011101011: begin rgb_reg = 3'b111; end
            18'b100000110011101100: begin rgb_reg = 3'b111; end
            18'b100000110011101101: begin rgb_reg = 3'b111; end
            18'b100000110011101110: begin rgb_reg = 3'b111; end
            18'b100000110011110110: begin rgb_reg = 3'b111; end
            18'b100000110011110111: begin rgb_reg = 3'b111; end
            18'b100000110011111000: begin rgb_reg = 3'b111; end
            18'b100000110011111001: begin rgb_reg = 3'b111; end
            18'b100000110011111010: begin rgb_reg = 3'b111; end
            18'b100000110011111011: begin rgb_reg = 3'b111; end
            18'b100000110011111100: begin rgb_reg = 3'b111; end
            18'b100000110100000011: begin rgb_reg = 3'b111; end
            18'b100000110100000100: begin rgb_reg = 3'b111; end
            18'b100000110100000101: begin rgb_reg = 3'b111; end
            18'b100000110100000110: begin rgb_reg = 3'b111; end
            18'b100000110100000111: begin rgb_reg = 3'b111; end
            18'b100000110100001000: begin rgb_reg = 3'b111; end
            18'b100000110100001001: begin rgb_reg = 3'b111; end
            18'b100000110100010011: begin rgb_reg = 3'b111; end
            18'b100000110100010100: begin rgb_reg = 3'b111; end
            18'b100000110100010101: begin rgb_reg = 3'b111; end
            18'b100000110100010110: begin rgb_reg = 3'b111; end
            18'b100000110100010111: begin rgb_reg = 3'b111; end
            18'b100000110100100001: begin rgb_reg = 3'b111; end
            18'b100000110100100010: begin rgb_reg = 3'b111; end
            18'b100000110100101100: begin rgb_reg = 3'b111; end
            18'b100000110100101101: begin rgb_reg = 3'b111; end
            18'b100000110100101110: begin rgb_reg = 3'b111; end
            18'b100000110100101111: begin rgb_reg = 3'b111; end
            18'b100000110100110000: begin rgb_reg = 3'b111; end
            18'b100000110100110001: begin rgb_reg = 3'b111; end
            18'b100000110100110010: begin rgb_reg = 3'b111; end
            18'b100000110100111100: begin rgb_reg = 3'b111; end
            18'b100000110100111101: begin rgb_reg = 3'b111; end
            18'b100000111011000000: begin rgb_reg = 3'b111; end
            18'b100000111011000001: begin rgb_reg = 3'b111; end
            18'b100000111011001011: begin rgb_reg = 3'b111; end
            18'b100000111011001100: begin rgb_reg = 3'b111; end
            18'b100000111011001101: begin rgb_reg = 3'b111; end
            18'b100000111011010100: begin rgb_reg = 3'b111; end
            18'b100000111011010101: begin rgb_reg = 3'b111; end
            18'b100000111011011001: begin rgb_reg = 3'b111; end
            18'b100000111011011010: begin rgb_reg = 3'b111; end
            18'b100000111011100010: begin rgb_reg = 3'b111; end
            18'b100000111011100011: begin rgb_reg = 3'b111; end
            18'b100000111011100110: begin rgb_reg = 3'b111; end
            18'b100000111011100111: begin rgb_reg = 3'b111; end
            18'b100000111011101000: begin rgb_reg = 3'b111; end
            18'b100000111011101111: begin rgb_reg = 3'b111; end
            18'b100000111011110000: begin rgb_reg = 3'b111; end
            18'b100000111011110100: begin rgb_reg = 3'b111; end
            18'b100000111011110101: begin rgb_reg = 3'b111; end
            18'b100000111011111101: begin rgb_reg = 3'b111; end
            18'b100000111011111110: begin rgb_reg = 3'b111; end
            18'b100000111100000001: begin rgb_reg = 3'b111; end
            18'b100000111100000010: begin rgb_reg = 3'b111; end
            18'b100000111100000011: begin rgb_reg = 3'b111; end
            18'b100000111100001010: begin rgb_reg = 3'b111; end
            18'b100000111100001011: begin rgb_reg = 3'b111; end
            18'b100000111100010001: begin rgb_reg = 3'b111; end
            18'b100000111100010010: begin rgb_reg = 3'b111; end
            18'b100000111100011111: begin rgb_reg = 3'b111; end
            18'b100000111100100000: begin rgb_reg = 3'b111; end
            18'b100000111100100001: begin rgb_reg = 3'b111; end
            18'b100000111100100010: begin rgb_reg = 3'b111; end
            18'b100000111100101010: begin rgb_reg = 3'b111; end
            18'b100000111100101011: begin rgb_reg = 3'b111; end
            18'b100000111100110011: begin rgb_reg = 3'b111; end
            18'b100000111100110100: begin rgb_reg = 3'b111; end
            18'b100000111100111010: begin rgb_reg = 3'b111; end
            18'b100000111100111011: begin rgb_reg = 3'b111; end
            18'b100000111100111100: begin rgb_reg = 3'b111; end
            18'b100000111100111101: begin rgb_reg = 3'b111; end
            18'b100001000011000000: begin rgb_reg = 3'b111; end
            18'b100001000011000001: begin rgb_reg = 3'b111; end
            18'b100001000011001011: begin rgb_reg = 3'b111; end
            18'b100001000011001100: begin rgb_reg = 3'b111; end
            18'b100001000011001101: begin rgb_reg = 3'b111; end
            18'b100001000011010100: begin rgb_reg = 3'b111; end
            18'b100001000011010101: begin rgb_reg = 3'b111; end
            18'b100001000011010110: begin rgb_reg = 3'b111; end
            18'b100001000011011001: begin rgb_reg = 3'b111; end
            18'b100001000011011010: begin rgb_reg = 3'b111; end
            18'b100001000011100010: begin rgb_reg = 3'b111; end
            18'b100001000011100011: begin rgb_reg = 3'b111; end
            18'b100001000011100110: begin rgb_reg = 3'b111; end
            18'b100001000011100111: begin rgb_reg = 3'b111; end
            18'b100001000011101000: begin rgb_reg = 3'b111; end
            18'b100001000011101111: begin rgb_reg = 3'b111; end
            18'b100001000011110000: begin rgb_reg = 3'b111; end
            18'b100001000011110001: begin rgb_reg = 3'b111; end
            18'b100001000011110100: begin rgb_reg = 3'b111; end
            18'b100001000011110101: begin rgb_reg = 3'b111; end
            18'b100001000011111101: begin rgb_reg = 3'b111; end
            18'b100001000011111110: begin rgb_reg = 3'b111; end
            18'b100001000100000001: begin rgb_reg = 3'b111; end
            18'b100001000100000010: begin rgb_reg = 3'b111; end
            18'b100001000100000011: begin rgb_reg = 3'b111; end
            18'b100001000100001010: begin rgb_reg = 3'b111; end
            18'b100001000100001011: begin rgb_reg = 3'b111; end
            18'b100001000100001100: begin rgb_reg = 3'b111; end
            18'b100001000100010001: begin rgb_reg = 3'b111; end
            18'b100001000100010010: begin rgb_reg = 3'b111; end
            18'b100001000100011110: begin rgb_reg = 3'b111; end
            18'b100001000100011111: begin rgb_reg = 3'b111; end
            18'b100001000100100000: begin rgb_reg = 3'b111; end
            18'b100001000100100001: begin rgb_reg = 3'b111; end
            18'b100001000100100010: begin rgb_reg = 3'b111; end
            18'b100001000100101010: begin rgb_reg = 3'b111; end
            18'b100001000100101011: begin rgb_reg = 3'b111; end
            18'b100001000100110011: begin rgb_reg = 3'b111; end
            18'b100001000100110100: begin rgb_reg = 3'b111; end
            18'b100001000100111001: begin rgb_reg = 3'b111; end
            18'b100001000100111010: begin rgb_reg = 3'b111; end
            18'b100001000100111011: begin rgb_reg = 3'b111; end
            18'b100001000100111100: begin rgb_reg = 3'b111; end
            18'b100001000100111101: begin rgb_reg = 3'b111; end
            18'b100001001010111110: begin rgb_reg = 3'b111; end
            18'b100001001010111111: begin rgb_reg = 3'b111; end
            18'b100001001011000000: begin rgb_reg = 3'b111; end
            18'b100001001011000001: begin rgb_reg = 3'b111; end
            18'b100001001011001011: begin rgb_reg = 3'b111; end
            18'b100001001011001100: begin rgb_reg = 3'b111; end
            18'b100001001011001101: begin rgb_reg = 3'b111; end
            18'b100001001011010010: begin rgb_reg = 3'b111; end
            18'b100001001011010011: begin rgb_reg = 3'b111; end
            18'b100001001011010100: begin rgb_reg = 3'b111; end
            18'b100001001011010101: begin rgb_reg = 3'b111; end
            18'b100001001011010110: begin rgb_reg = 3'b111; end
            18'b100001001011011001: begin rgb_reg = 3'b111; end
            18'b100001001011011010: begin rgb_reg = 3'b111; end
            18'b100001001011100010: begin rgb_reg = 3'b111; end
            18'b100001001011100011: begin rgb_reg = 3'b111; end
            18'b100001001011100110: begin rgb_reg = 3'b111; end
            18'b100001001011100111: begin rgb_reg = 3'b111; end
            18'b100001001011101000: begin rgb_reg = 3'b111; end
            18'b100001001011101101: begin rgb_reg = 3'b111; end
            18'b100001001011101110: begin rgb_reg = 3'b111; end
            18'b100001001011101111: begin rgb_reg = 3'b111; end
            18'b100001001011110000: begin rgb_reg = 3'b111; end
            18'b100001001011110001: begin rgb_reg = 3'b111; end
            18'b100001001011110100: begin rgb_reg = 3'b111; end
            18'b100001001011110101: begin rgb_reg = 3'b111; end
            18'b100001001011111101: begin rgb_reg = 3'b111; end
            18'b100001001011111110: begin rgb_reg = 3'b111; end
            18'b100001001100000010: begin rgb_reg = 3'b111; end
            18'b100001001100001010: begin rgb_reg = 3'b111; end
            18'b100001001100001011: begin rgb_reg = 3'b111; end
            18'b100001001100001100: begin rgb_reg = 3'b111; end
            18'b100001001100001111: begin rgb_reg = 3'b111; end
            18'b100001001100010000: begin rgb_reg = 3'b111; end
            18'b100001001100010001: begin rgb_reg = 3'b111; end
            18'b100001001100010010: begin rgb_reg = 3'b111; end
            18'b100001001100011111: begin rgb_reg = 3'b111; end
            18'b100001001100100000: begin rgb_reg = 3'b111; end
            18'b100001001100100001: begin rgb_reg = 3'b111; end
            18'b100001001100100010: begin rgb_reg = 3'b111; end
            18'b100001001100101010: begin rgb_reg = 3'b111; end
            18'b100001001100101011: begin rgb_reg = 3'b111; end
            18'b100001001100110011: begin rgb_reg = 3'b111; end
            18'b100001001100110100: begin rgb_reg = 3'b111; end
            18'b100001001100111010: begin rgb_reg = 3'b111; end
            18'b100001001100111011: begin rgb_reg = 3'b111; end
            18'b100001001100111100: begin rgb_reg = 3'b111; end
            18'b100001001100111101: begin rgb_reg = 3'b111; end
            18'b100001010010111110: begin rgb_reg = 3'b111; end
            18'b100001010010111111: begin rgb_reg = 3'b111; end
            18'b100001010011001011: begin rgb_reg = 3'b111; end
            18'b100001010011001100: begin rgb_reg = 3'b111; end
            18'b100001010011001101: begin rgb_reg = 3'b111; end
            18'b100001010011010010: begin rgb_reg = 3'b111; end
            18'b100001010011010011: begin rgb_reg = 3'b111; end
            18'b100001010011010100: begin rgb_reg = 3'b111; end
            18'b100001010011010101: begin rgb_reg = 3'b111; end
            18'b100001010011010110: begin rgb_reg = 3'b111; end
            18'b100001010011100010: begin rgb_reg = 3'b111; end
            18'b100001010011100011: begin rgb_reg = 3'b111; end
            18'b100001010011100110: begin rgb_reg = 3'b111; end
            18'b100001010011100111: begin rgb_reg = 3'b111; end
            18'b100001010011101000: begin rgb_reg = 3'b111; end
            18'b100001010011101101: begin rgb_reg = 3'b111; end
            18'b100001010011101110: begin rgb_reg = 3'b111; end
            18'b100001010011101111: begin rgb_reg = 3'b111; end
            18'b100001010011110000: begin rgb_reg = 3'b111; end
            18'b100001010011110001: begin rgb_reg = 3'b111; end
            18'b100001010011111101: begin rgb_reg = 3'b111; end
            18'b100001010011111110: begin rgb_reg = 3'b111; end
            18'b100001010100001010: begin rgb_reg = 3'b111; end
            18'b100001010100001011: begin rgb_reg = 3'b111; end
            18'b100001010100001100: begin rgb_reg = 3'b111; end
            18'b100001010100001111: begin rgb_reg = 3'b111; end
            18'b100001010100010000: begin rgb_reg = 3'b111; end
            18'b100001010100100001: begin rgb_reg = 3'b111; end
            18'b100001010100100010: begin rgb_reg = 3'b111; end
            18'b100001010100110011: begin rgb_reg = 3'b111; end
            18'b100001010100110100: begin rgb_reg = 3'b111; end
            18'b100001010100111100: begin rgb_reg = 3'b111; end
            18'b100001010100111101: begin rgb_reg = 3'b111; end
            18'b100001011010111110: begin rgb_reg = 3'b111; end
            18'b100001011010111111: begin rgb_reg = 3'b111; end
            18'b100001011011001011: begin rgb_reg = 3'b111; end
            18'b100001011011001100: begin rgb_reg = 3'b111; end
            18'b100001011011001101: begin rgb_reg = 3'b111; end
            18'b100001011011010010: begin rgb_reg = 3'b111; end
            18'b100001011011010011: begin rgb_reg = 3'b111; end
            18'b100001011011010100: begin rgb_reg = 3'b111; end
            18'b100001011011010101: begin rgb_reg = 3'b111; end
            18'b100001011011010110: begin rgb_reg = 3'b111; end
            18'b100001011011100010: begin rgb_reg = 3'b111; end
            18'b100001011011100011: begin rgb_reg = 3'b111; end
            18'b100001011011100110: begin rgb_reg = 3'b111; end
            18'b100001011011100111: begin rgb_reg = 3'b111; end
            18'b100001011011101000: begin rgb_reg = 3'b111; end
            18'b100001011011101101: begin rgb_reg = 3'b111; end
            18'b100001011011101110: begin rgb_reg = 3'b111; end
            18'b100001011011101111: begin rgb_reg = 3'b111; end
            18'b100001011011110000: begin rgb_reg = 3'b111; end
            18'b100001011011110001: begin rgb_reg = 3'b111; end
            18'b100001011011111101: begin rgb_reg = 3'b111; end
            18'b100001011011111110: begin rgb_reg = 3'b111; end
            18'b100001011100001010: begin rgb_reg = 3'b111; end
            18'b100001011100001011: begin rgb_reg = 3'b111; end
            18'b100001011100001111: begin rgb_reg = 3'b111; end
            18'b100001011100010000: begin rgb_reg = 3'b111; end
            18'b100001011100100001: begin rgb_reg = 3'b111; end
            18'b100001011100100010: begin rgb_reg = 3'b111; end
            18'b100001011100110011: begin rgb_reg = 3'b111; end
            18'b100001011100110100: begin rgb_reg = 3'b111; end
            18'b100001011100111100: begin rgb_reg = 3'b111; end
            18'b100001011100111101: begin rgb_reg = 3'b111; end
            18'b100001100010111110: begin rgb_reg = 3'b111; end
            18'b100001100010111111: begin rgb_reg = 3'b111; end
            18'b100001100011000000: begin rgb_reg = 3'b111; end
            18'b100001100011000001: begin rgb_reg = 3'b111; end
            18'b100001100011000010: begin rgb_reg = 3'b111; end
            18'b100001100011000011: begin rgb_reg = 3'b111; end
            18'b100001100011000100: begin rgb_reg = 3'b111; end
            18'b100001100011000101: begin rgb_reg = 3'b111; end
            18'b100001100011000110: begin rgb_reg = 3'b111; end
            18'b100001100011001011: begin rgb_reg = 3'b111; end
            18'b100001100011001100: begin rgb_reg = 3'b111; end
            18'b100001100011001101: begin rgb_reg = 3'b111; end
            18'b100001100011010000: begin rgb_reg = 3'b111; end
            18'b100001100011010001: begin rgb_reg = 3'b111; end
            18'b100001100011010100: begin rgb_reg = 3'b111; end
            18'b100001100011010101: begin rgb_reg = 3'b111; end
            18'b100001100011010110: begin rgb_reg = 3'b111; end
            18'b100001100011011101: begin rgb_reg = 3'b111; end
            18'b100001100011011110: begin rgb_reg = 3'b111; end
            18'b100001100011011111: begin rgb_reg = 3'b111; end
            18'b100001100011100000: begin rgb_reg = 3'b111; end
            18'b100001100011100001: begin rgb_reg = 3'b111; end
            18'b100001100011100110: begin rgb_reg = 3'b111; end
            18'b100001100011100111: begin rgb_reg = 3'b111; end
            18'b100001100011101000: begin rgb_reg = 3'b111; end
            18'b100001100011101011: begin rgb_reg = 3'b111; end
            18'b100001100011101100: begin rgb_reg = 3'b111; end
            18'b100001100011101111: begin rgb_reg = 3'b111; end
            18'b100001100011110000: begin rgb_reg = 3'b111; end
            18'b100001100011110001: begin rgb_reg = 3'b111; end
            18'b100001100011111000: begin rgb_reg = 3'b111; end
            18'b100001100011111001: begin rgb_reg = 3'b111; end
            18'b100001100011111010: begin rgb_reg = 3'b111; end
            18'b100001100011111011: begin rgb_reg = 3'b111; end
            18'b100001100011111100: begin rgb_reg = 3'b111; end
            18'b100001100100000110: begin rgb_reg = 3'b111; end
            18'b100001100100000111: begin rgb_reg = 3'b111; end
            18'b100001100100001000: begin rgb_reg = 3'b111; end
            18'b100001100100001001: begin rgb_reg = 3'b111; end
            18'b100001100100001111: begin rgb_reg = 3'b111; end
            18'b100001100100010000: begin rgb_reg = 3'b111; end
            18'b100001100100010001: begin rgb_reg = 3'b111; end
            18'b100001100100010010: begin rgb_reg = 3'b111; end
            18'b100001100100010011: begin rgb_reg = 3'b111; end
            18'b100001100100010100: begin rgb_reg = 3'b111; end
            18'b100001100100010101: begin rgb_reg = 3'b111; end
            18'b100001100100010110: begin rgb_reg = 3'b111; end
            18'b100001100100010111: begin rgb_reg = 3'b111; end
            18'b100001100100100001: begin rgb_reg = 3'b111; end
            18'b100001100100100010: begin rgb_reg = 3'b111; end
            18'b100001100100101110: begin rgb_reg = 3'b111; end
            18'b100001100100101111: begin rgb_reg = 3'b111; end
            18'b100001100100110000: begin rgb_reg = 3'b111; end
            18'b100001100100110001: begin rgb_reg = 3'b111; end
            18'b100001100100110010: begin rgb_reg = 3'b111; end
            18'b100001100100111100: begin rgb_reg = 3'b111; end
            18'b100001100100111101: begin rgb_reg = 3'b111; end
            18'b100001101010111110: begin rgb_reg = 3'b111; end
            18'b100001101010111111: begin rgb_reg = 3'b111; end
            18'b100001101011000000: begin rgb_reg = 3'b111; end
            18'b100001101011000001: begin rgb_reg = 3'b111; end
            18'b100001101011000010: begin rgb_reg = 3'b111; end
            18'b100001101011000011: begin rgb_reg = 3'b111; end
            18'b100001101011000100: begin rgb_reg = 3'b111; end
            18'b100001101011000101: begin rgb_reg = 3'b111; end
            18'b100001101011000110: begin rgb_reg = 3'b111; end
            18'b100001101011001011: begin rgb_reg = 3'b111; end
            18'b100001101011001100: begin rgb_reg = 3'b111; end
            18'b100001101011001101: begin rgb_reg = 3'b111; end
            18'b100001101011010000: begin rgb_reg = 3'b111; end
            18'b100001101011010001: begin rgb_reg = 3'b111; end
            18'b100001101011010100: begin rgb_reg = 3'b111; end
            18'b100001101011010101: begin rgb_reg = 3'b111; end
            18'b100001101011010110: begin rgb_reg = 3'b111; end
            18'b100001101011011101: begin rgb_reg = 3'b111; end
            18'b100001101011011110: begin rgb_reg = 3'b111; end
            18'b100001101011011111: begin rgb_reg = 3'b111; end
            18'b100001101011100000: begin rgb_reg = 3'b111; end
            18'b100001101011100001: begin rgb_reg = 3'b111; end
            18'b100001101011100110: begin rgb_reg = 3'b111; end
            18'b100001101011100111: begin rgb_reg = 3'b111; end
            18'b100001101011101000: begin rgb_reg = 3'b111; end
            18'b100001101011101011: begin rgb_reg = 3'b111; end
            18'b100001101011101100: begin rgb_reg = 3'b111; end
            18'b100001101011101111: begin rgb_reg = 3'b111; end
            18'b100001101011110000: begin rgb_reg = 3'b111; end
            18'b100001101011110001: begin rgb_reg = 3'b111; end
            18'b100001101011111000: begin rgb_reg = 3'b111; end
            18'b100001101011111001: begin rgb_reg = 3'b111; end
            18'b100001101011111010: begin rgb_reg = 3'b111; end
            18'b100001101011111011: begin rgb_reg = 3'b111; end
            18'b100001101011111100: begin rgb_reg = 3'b111; end
            18'b100001101100000110: begin rgb_reg = 3'b111; end
            18'b100001101100000111: begin rgb_reg = 3'b111; end
            18'b100001101100001000: begin rgb_reg = 3'b111; end
            18'b100001101100001001: begin rgb_reg = 3'b111; end
            18'b100001101100001111: begin rgb_reg = 3'b111; end
            18'b100001101100010000: begin rgb_reg = 3'b111; end
            18'b100001101100010001: begin rgb_reg = 3'b111; end
            18'b100001101100010010: begin rgb_reg = 3'b111; end
            18'b100001101100010011: begin rgb_reg = 3'b111; end
            18'b100001101100010100: begin rgb_reg = 3'b111; end
            18'b100001101100010101: begin rgb_reg = 3'b111; end
            18'b100001101100010110: begin rgb_reg = 3'b111; end
            18'b100001101100010111: begin rgb_reg = 3'b111; end
            18'b100001101100100001: begin rgb_reg = 3'b111; end
            18'b100001101100100010: begin rgb_reg = 3'b111; end
            18'b100001101100101110: begin rgb_reg = 3'b111; end
            18'b100001101100101111: begin rgb_reg = 3'b111; end
            18'b100001101100110000: begin rgb_reg = 3'b111; end
            18'b100001101100110001: begin rgb_reg = 3'b111; end
            18'b100001101100110010: begin rgb_reg = 3'b111; end
            18'b100001101100111100: begin rgb_reg = 3'b111; end
            18'b100001101100111101: begin rgb_reg = 3'b111; end
            18'b100001110010111110: begin rgb_reg = 3'b111; end
            18'b100001110010111111: begin rgb_reg = 3'b111; end
            18'b100001110011000111: begin rgb_reg = 3'b111; end
            18'b100001110011001000: begin rgb_reg = 3'b111; end
            18'b100001110011001011: begin rgb_reg = 3'b111; end
            18'b100001110011001100: begin rgb_reg = 3'b111; end
            18'b100001110011001101: begin rgb_reg = 3'b111; end
            18'b100001110011001110: begin rgb_reg = 3'b111; end
            18'b100001110011001111: begin rgb_reg = 3'b111; end
            18'b100001110011010100: begin rgb_reg = 3'b111; end
            18'b100001110011010101: begin rgb_reg = 3'b111; end
            18'b100001110011010110: begin rgb_reg = 3'b111; end
            18'b100001110011100010: begin rgb_reg = 3'b111; end
            18'b100001110011100011: begin rgb_reg = 3'b111; end
            18'b100001110011100110: begin rgb_reg = 3'b111; end
            18'b100001110011100111: begin rgb_reg = 3'b111; end
            18'b100001110011101000: begin rgb_reg = 3'b111; end
            18'b100001110011101001: begin rgb_reg = 3'b111; end
            18'b100001110011101010: begin rgb_reg = 3'b111; end
            18'b100001110011101111: begin rgb_reg = 3'b111; end
            18'b100001110011110000: begin rgb_reg = 3'b111; end
            18'b100001110011110001: begin rgb_reg = 3'b111; end
            18'b100001110011110110: begin rgb_reg = 3'b111; end
            18'b100001110011110111: begin rgb_reg = 3'b111; end
            18'b100001110100000011: begin rgb_reg = 3'b111; end
            18'b100001110100000100: begin rgb_reg = 3'b111; end
            18'b100001110100000101: begin rgb_reg = 3'b111; end
            18'b100001110100001111: begin rgb_reg = 3'b111; end
            18'b100001110100010000: begin rgb_reg = 3'b111; end
            18'b100001110100011000: begin rgb_reg = 3'b111; end
            18'b100001110100011001: begin rgb_reg = 3'b111; end
            18'b100001110100100001: begin rgb_reg = 3'b111; end
            18'b100001110100100010: begin rgb_reg = 3'b111; end
            18'b100001110100101100: begin rgb_reg = 3'b111; end
            18'b100001110100101101: begin rgb_reg = 3'b111; end
            18'b100001110100111100: begin rgb_reg = 3'b111; end
            18'b100001110100111101: begin rgb_reg = 3'b111; end
            18'b100001111010111110: begin rgb_reg = 3'b111; end
            18'b100001111010111111: begin rgb_reg = 3'b111; end
            18'b100001111011000111: begin rgb_reg = 3'b111; end
            18'b100001111011001000: begin rgb_reg = 3'b111; end
            18'b100001111011001011: begin rgb_reg = 3'b111; end
            18'b100001111011001100: begin rgb_reg = 3'b111; end
            18'b100001111011001101: begin rgb_reg = 3'b111; end
            18'b100001111011001110: begin rgb_reg = 3'b111; end
            18'b100001111011001111: begin rgb_reg = 3'b111; end
            18'b100001111011010100: begin rgb_reg = 3'b111; end
            18'b100001111011010101: begin rgb_reg = 3'b111; end
            18'b100001111011010110: begin rgb_reg = 3'b111; end
            18'b100001111011100010: begin rgb_reg = 3'b111; end
            18'b100001111011100011: begin rgb_reg = 3'b111; end
            18'b100001111011100110: begin rgb_reg = 3'b111; end
            18'b100001111011100111: begin rgb_reg = 3'b111; end
            18'b100001111011101000: begin rgb_reg = 3'b111; end
            18'b100001111011101001: begin rgb_reg = 3'b111; end
            18'b100001111011101010: begin rgb_reg = 3'b111; end
            18'b100001111011101111: begin rgb_reg = 3'b111; end
            18'b100001111011110000: begin rgb_reg = 3'b111; end
            18'b100001111011110001: begin rgb_reg = 3'b111; end
            18'b100001111011110110: begin rgb_reg = 3'b111; end
            18'b100001111011110111: begin rgb_reg = 3'b111; end
            18'b100001111100000011: begin rgb_reg = 3'b111; end
            18'b100001111100000100: begin rgb_reg = 3'b111; end
            18'b100001111100000101: begin rgb_reg = 3'b111; end
            18'b100001111100001111: begin rgb_reg = 3'b111; end
            18'b100001111100010000: begin rgb_reg = 3'b111; end
            18'b100001111100011000: begin rgb_reg = 3'b111; end
            18'b100001111100011001: begin rgb_reg = 3'b111; end
            18'b100001111100100001: begin rgb_reg = 3'b111; end
            18'b100001111100100010: begin rgb_reg = 3'b111; end
            18'b100001111100101100: begin rgb_reg = 3'b111; end
            18'b100001111100101101: begin rgb_reg = 3'b111; end
            18'b100001111100111100: begin rgb_reg = 3'b111; end
            18'b100001111100111101: begin rgb_reg = 3'b111; end
            18'b100010000010111110: begin rgb_reg = 3'b111; end
            18'b100010000010111111: begin rgb_reg = 3'b111; end
            18'b100010000011000111: begin rgb_reg = 3'b111; end
            18'b100010000011001000: begin rgb_reg = 3'b111; end
            18'b100010000011001011: begin rgb_reg = 3'b111; end
            18'b100010000011001100: begin rgb_reg = 3'b111; end
            18'b100010000011001101: begin rgb_reg = 3'b111; end
            18'b100010000011010100: begin rgb_reg = 3'b111; end
            18'b100010000011010101: begin rgb_reg = 3'b111; end
            18'b100010000011010110: begin rgb_reg = 3'b111; end
            18'b100010000011011001: begin rgb_reg = 3'b111; end
            18'b100010000011011010: begin rgb_reg = 3'b111; end
            18'b100010000011100010: begin rgb_reg = 3'b111; end
            18'b100010000011100011: begin rgb_reg = 3'b111; end
            18'b100010000011100110: begin rgb_reg = 3'b111; end
            18'b100010000011100111: begin rgb_reg = 3'b111; end
            18'b100010000011101000: begin rgb_reg = 3'b111; end
            18'b100010000011101111: begin rgb_reg = 3'b111; end
            18'b100010000011110000: begin rgb_reg = 3'b111; end
            18'b100010000011110001: begin rgb_reg = 3'b111; end
            18'b100010000011110100: begin rgb_reg = 3'b111; end
            18'b100010000011110101: begin rgb_reg = 3'b111; end
            18'b100010000100000001: begin rgb_reg = 3'b111; end
            18'b100010000100000010: begin rgb_reg = 3'b111; end
            18'b100010000100000011: begin rgb_reg = 3'b111; end
            18'b100010000100001111: begin rgb_reg = 3'b111; end
            18'b100010000100010000: begin rgb_reg = 3'b111; end
            18'b100010000100011000: begin rgb_reg = 3'b111; end
            18'b100010000100011001: begin rgb_reg = 3'b111; end
            18'b100010000100100001: begin rgb_reg = 3'b111; end
            18'b100010000100100010: begin rgb_reg = 3'b111; end
            18'b100010000100101010: begin rgb_reg = 3'b111; end
            18'b100010000100101011: begin rgb_reg = 3'b111; end
            18'b100010000100111100: begin rgb_reg = 3'b111; end
            18'b100010000100111101: begin rgb_reg = 3'b111; end
            18'b100010001010111110: begin rgb_reg = 3'b111; end
            18'b100010001010111111: begin rgb_reg = 3'b111; end
            18'b100010001011000111: begin rgb_reg = 3'b111; end
            18'b100010001011001000: begin rgb_reg = 3'b111; end
            18'b100010001011001011: begin rgb_reg = 3'b111; end
            18'b100010001011001100: begin rgb_reg = 3'b111; end
            18'b100010001011001101: begin rgb_reg = 3'b111; end
            18'b100010001011010100: begin rgb_reg = 3'b111; end
            18'b100010001011010101: begin rgb_reg = 3'b111; end
            18'b100010001011010110: begin rgb_reg = 3'b111; end
            18'b100010001011011001: begin rgb_reg = 3'b111; end
            18'b100010001011011010: begin rgb_reg = 3'b111; end
            18'b100010001011100010: begin rgb_reg = 3'b111; end
            18'b100010001011100011: begin rgb_reg = 3'b111; end
            18'b100010001011100110: begin rgb_reg = 3'b111; end
            18'b100010001011100111: begin rgb_reg = 3'b111; end
            18'b100010001011101000: begin rgb_reg = 3'b111; end
            18'b100010001011101111: begin rgb_reg = 3'b111; end
            18'b100010001011110000: begin rgb_reg = 3'b111; end
            18'b100010001011110001: begin rgb_reg = 3'b111; end
            18'b100010001011110100: begin rgb_reg = 3'b111; end
            18'b100010001011110101: begin rgb_reg = 3'b111; end
            18'b100010001100000001: begin rgb_reg = 3'b111; end
            18'b100010001100000010: begin rgb_reg = 3'b111; end
            18'b100010001100000011: begin rgb_reg = 3'b111; end
            18'b100010001100001111: begin rgb_reg = 3'b111; end
            18'b100010001100010000: begin rgb_reg = 3'b111; end
            18'b100010001100011000: begin rgb_reg = 3'b111; end
            18'b100010001100011001: begin rgb_reg = 3'b111; end
            18'b100010001100100001: begin rgb_reg = 3'b111; end
            18'b100010001100100010: begin rgb_reg = 3'b111; end
            18'b100010001100101010: begin rgb_reg = 3'b111; end
            18'b100010001100101011: begin rgb_reg = 3'b111; end
            18'b100010001100111100: begin rgb_reg = 3'b111; end
            18'b100010001100111101: begin rgb_reg = 3'b111; end
            18'b100010010010111110: begin rgb_reg = 3'b111; end
            18'b100010010010111111: begin rgb_reg = 3'b111; end
            18'b100010010011000000: begin rgb_reg = 3'b111; end
            18'b100010010011000001: begin rgb_reg = 3'b111; end
            18'b100010010011000010: begin rgb_reg = 3'b111; end
            18'b100010010011000011: begin rgb_reg = 3'b111; end
            18'b100010010011000100: begin rgb_reg = 3'b111; end
            18'b100010010011000101: begin rgb_reg = 3'b111; end
            18'b100010010011000110: begin rgb_reg = 3'b111; end
            18'b100010010011000111: begin rgb_reg = 3'b111; end
            18'b100010010011001000: begin rgb_reg = 3'b111; end
            18'b100010010011001100: begin rgb_reg = 3'b111; end
            18'b100010010011001101: begin rgb_reg = 3'b111; end
            18'b100010010011001110: begin rgb_reg = 3'b111; end
            18'b100010010011001111: begin rgb_reg = 3'b111; end
            18'b100010010011010000: begin rgb_reg = 3'b111; end
            18'b100010010011010001: begin rgb_reg = 3'b111; end
            18'b100010010011010010: begin rgb_reg = 3'b111; end
            18'b100010010011010011: begin rgb_reg = 3'b111; end
            18'b100010010011010100: begin rgb_reg = 3'b111; end
            18'b100010010011010101: begin rgb_reg = 3'b111; end
            18'b100010010011011001: begin rgb_reg = 3'b111; end
            18'b100010010011011010: begin rgb_reg = 3'b111; end
            18'b100010010011011011: begin rgb_reg = 3'b111; end
            18'b100010010011011100: begin rgb_reg = 3'b111; end
            18'b100010010011011101: begin rgb_reg = 3'b111; end
            18'b100010010011011110: begin rgb_reg = 3'b111; end
            18'b100010010011011111: begin rgb_reg = 3'b111; end
            18'b100010010011100000: begin rgb_reg = 3'b111; end
            18'b100010010011100001: begin rgb_reg = 3'b111; end
            18'b100010010011100010: begin rgb_reg = 3'b111; end
            18'b100010010011100011: begin rgb_reg = 3'b111; end
            18'b100010010011100111: begin rgb_reg = 3'b111; end
            18'b100010010011101000: begin rgb_reg = 3'b111; end
            18'b100010010011101001: begin rgb_reg = 3'b111; end
            18'b100010010011101010: begin rgb_reg = 3'b111; end
            18'b100010010011101011: begin rgb_reg = 3'b111; end
            18'b100010010011101100: begin rgb_reg = 3'b111; end
            18'b100010010011101101: begin rgb_reg = 3'b111; end
            18'b100010010011101110: begin rgb_reg = 3'b111; end
            18'b100010010011101111: begin rgb_reg = 3'b111; end
            18'b100010010011110000: begin rgb_reg = 3'b111; end
            18'b100010010011110100: begin rgb_reg = 3'b111; end
            18'b100010010011110101: begin rgb_reg = 3'b111; end
            18'b100010010011110110: begin rgb_reg = 3'b111; end
            18'b100010010011110111: begin rgb_reg = 3'b111; end
            18'b100010010011111000: begin rgb_reg = 3'b111; end
            18'b100010010011111001: begin rgb_reg = 3'b111; end
            18'b100010010011111010: begin rgb_reg = 3'b111; end
            18'b100010010011111011: begin rgb_reg = 3'b111; end
            18'b100010010011111100: begin rgb_reg = 3'b111; end
            18'b100010010011111101: begin rgb_reg = 3'b111; end
            18'b100010010011111110: begin rgb_reg = 3'b111; end
            18'b100010010100000001: begin rgb_reg = 3'b111; end
            18'b100010010100000010: begin rgb_reg = 3'b111; end
            18'b100010010100000011: begin rgb_reg = 3'b111; end
            18'b100010010100000100: begin rgb_reg = 3'b111; end
            18'b100010010100000101: begin rgb_reg = 3'b111; end
            18'b100010010100000110: begin rgb_reg = 3'b111; end
            18'b100010010100000111: begin rgb_reg = 3'b111; end
            18'b100010010100001000: begin rgb_reg = 3'b111; end
            18'b100010010100001001: begin rgb_reg = 3'b111; end
            18'b100010010100001010: begin rgb_reg = 3'b111; end
            18'b100010010100001011: begin rgb_reg = 3'b111; end
            18'b100010010100001111: begin rgb_reg = 3'b111; end
            18'b100010010100010000: begin rgb_reg = 3'b111; end
            18'b100010010100010001: begin rgb_reg = 3'b111; end
            18'b100010010100010010: begin rgb_reg = 3'b111; end
            18'b100010010100010011: begin rgb_reg = 3'b111; end
            18'b100010010100010100: begin rgb_reg = 3'b111; end
            18'b100010010100010101: begin rgb_reg = 3'b111; end
            18'b100010010100010110: begin rgb_reg = 3'b111; end
            18'b100010010100010111: begin rgb_reg = 3'b111; end
            18'b100010010100011000: begin rgb_reg = 3'b111; end
            18'b100010010100011001: begin rgb_reg = 3'b111; end
            18'b100010010100011101: begin rgb_reg = 3'b111; end
            18'b100010010100011110: begin rgb_reg = 3'b111; end
            18'b100010010100011111: begin rgb_reg = 3'b111; end
            18'b100010010100100000: begin rgb_reg = 3'b111; end
            18'b100010010100100001: begin rgb_reg = 3'b111; end
            18'b100010010100100010: begin rgb_reg = 3'b111; end
            18'b100010010100100011: begin rgb_reg = 3'b111; end
            18'b100010010100100100: begin rgb_reg = 3'b111; end
            18'b100010010100100101: begin rgb_reg = 3'b111; end
            18'b100010010100100110: begin rgb_reg = 3'b111; end
            18'b100010010100101010: begin rgb_reg = 3'b111; end
            18'b100010010100101011: begin rgb_reg = 3'b111; end
            18'b100010010100101100: begin rgb_reg = 3'b111; end
            18'b100010010100101101: begin rgb_reg = 3'b111; end
            18'b100010010100101110: begin rgb_reg = 3'b111; end
            18'b100010010100101111: begin rgb_reg = 3'b111; end
            18'b100010010100110000: begin rgb_reg = 3'b111; end
            18'b100010010100110001: begin rgb_reg = 3'b111; end
            18'b100010010100110010: begin rgb_reg = 3'b111; end
            18'b100010010100110011: begin rgb_reg = 3'b111; end
            18'b100010010100110100: begin rgb_reg = 3'b111; end
            18'b100010010100111000: begin rgb_reg = 3'b111; end
            18'b100010010100111001: begin rgb_reg = 3'b111; end
            18'b100010010100111010: begin rgb_reg = 3'b111; end
            18'b100010010100111011: begin rgb_reg = 3'b111; end
            18'b100010010100111100: begin rgb_reg = 3'b111; end
            18'b100010010100111101: begin rgb_reg = 3'b111; end
            18'b100010010100111110: begin rgb_reg = 3'b111; end
            18'b100010010100111111: begin rgb_reg = 3'b111; end
            18'b100010010101000000: begin rgb_reg = 3'b111; end
            18'b100010010101000001: begin rgb_reg = 3'b111; end
            18'b100010011011000000: begin rgb_reg = 3'b111; end
            18'b100010011011000001: begin rgb_reg = 3'b111; end
            18'b100010011011000010: begin rgb_reg = 3'b111; end
            18'b100010011011000011: begin rgb_reg = 3'b111; end
            18'b100010011011000100: begin rgb_reg = 3'b111; end
            18'b100010011011000101: begin rgb_reg = 3'b111; end
            18'b100010011011000110: begin rgb_reg = 3'b111; end
            18'b100010011011001101: begin rgb_reg = 3'b111; end
            18'b100010011011001110: begin rgb_reg = 3'b111; end
            18'b100010011011001111: begin rgb_reg = 3'b111; end
            18'b100010011011010000: begin rgb_reg = 3'b111; end
            18'b100010011011010001: begin rgb_reg = 3'b111; end
            18'b100010011011010010: begin rgb_reg = 3'b111; end
            18'b100010011011010011: begin rgb_reg = 3'b111; end
            18'b100010011011011011: begin rgb_reg = 3'b111; end
            18'b100010011011011100: begin rgb_reg = 3'b111; end
            18'b100010011011011101: begin rgb_reg = 3'b111; end
            18'b100010011011011110: begin rgb_reg = 3'b111; end
            18'b100010011011011111: begin rgb_reg = 3'b111; end
            18'b100010011011100000: begin rgb_reg = 3'b111; end
            18'b100010011011100001: begin rgb_reg = 3'b111; end
            18'b100010011011101000: begin rgb_reg = 3'b111; end
            18'b100010011011101001: begin rgb_reg = 3'b111; end
            18'b100010011011101010: begin rgb_reg = 3'b111; end
            18'b100010011011101011: begin rgb_reg = 3'b111; end
            18'b100010011011101100: begin rgb_reg = 3'b111; end
            18'b100010011011101101: begin rgb_reg = 3'b111; end
            18'b100010011011101110: begin rgb_reg = 3'b111; end
            18'b100010011011110100: begin rgb_reg = 3'b111; end
            18'b100010011011110101: begin rgb_reg = 3'b111; end
            18'b100010011011110110: begin rgb_reg = 3'b111; end
            18'b100010011011110111: begin rgb_reg = 3'b111; end
            18'b100010011011111000: begin rgb_reg = 3'b111; end
            18'b100010011011111001: begin rgb_reg = 3'b111; end
            18'b100010011011111010: begin rgb_reg = 3'b111; end
            18'b100010011011111011: begin rgb_reg = 3'b111; end
            18'b100010011011111100: begin rgb_reg = 3'b111; end
            18'b100010011011111101: begin rgb_reg = 3'b111; end
            18'b100010011011111110: begin rgb_reg = 3'b111; end
            18'b100010011100000001: begin rgb_reg = 3'b111; end
            18'b100010011100000010: begin rgb_reg = 3'b111; end
            18'b100010011100000011: begin rgb_reg = 3'b111; end
            18'b100010011100000100: begin rgb_reg = 3'b111; end
            18'b100010011100000101: begin rgb_reg = 3'b111; end
            18'b100010011100000110: begin rgb_reg = 3'b111; end
            18'b100010011100000111: begin rgb_reg = 3'b111; end
            18'b100010011100001000: begin rgb_reg = 3'b111; end
            18'b100010011100001001: begin rgb_reg = 3'b111; end
            18'b100010011100001010: begin rgb_reg = 3'b111; end
            18'b100010011100001011: begin rgb_reg = 3'b111; end
            18'b100010011100001100: begin rgb_reg = 3'b111; end
            18'b100010011100010001: begin rgb_reg = 3'b111; end
            18'b100010011100010010: begin rgb_reg = 3'b111; end
            18'b100010011100010011: begin rgb_reg = 3'b111; end
            18'b100010011100010100: begin rgb_reg = 3'b111; end
            18'b100010011100010101: begin rgb_reg = 3'b111; end
            18'b100010011100010110: begin rgb_reg = 3'b111; end
            18'b100010011100010111: begin rgb_reg = 3'b111; end
            18'b100010011100011100: begin rgb_reg = 3'b111; end
            18'b100010011100011101: begin rgb_reg = 3'b111; end
            18'b100010011100011110: begin rgb_reg = 3'b111; end
            18'b100010011100011111: begin rgb_reg = 3'b111; end
            18'b100010011100100000: begin rgb_reg = 3'b111; end
            18'b100010011100100001: begin rgb_reg = 3'b111; end
            18'b100010011100100010: begin rgb_reg = 3'b111; end
            18'b100010011100100011: begin rgb_reg = 3'b111; end
            18'b100010011100100100: begin rgb_reg = 3'b111; end
            18'b100010011100100101: begin rgb_reg = 3'b111; end
            18'b100010011100100110: begin rgb_reg = 3'b111; end
            18'b100010011100100111: begin rgb_reg = 3'b111; end
            18'b100010011100101010: begin rgb_reg = 3'b111; end
            18'b100010011100101011: begin rgb_reg = 3'b111; end
            18'b100010011100101100: begin rgb_reg = 3'b111; end
            18'b100010011100101101: begin rgb_reg = 3'b111; end
            18'b100010011100101110: begin rgb_reg = 3'b111; end
            18'b100010011100101111: begin rgb_reg = 3'b111; end
            18'b100010011100110000: begin rgb_reg = 3'b111; end
            18'b100010011100110001: begin rgb_reg = 3'b111; end
            18'b100010011100110010: begin rgb_reg = 3'b111; end
            18'b100010011100110011: begin rgb_reg = 3'b111; end
            18'b100010011100110100: begin rgb_reg = 3'b111; end
            18'b100010011100110111: begin rgb_reg = 3'b111; end
            18'b100010011100111000: begin rgb_reg = 3'b111; end
            18'b100010011100111001: begin rgb_reg = 3'b111; end
            18'b100010011100111010: begin rgb_reg = 3'b111; end
            18'b100010011100111011: begin rgb_reg = 3'b111; end
            18'b100010011100111100: begin rgb_reg = 3'b111; end
            18'b100010011100111101: begin rgb_reg = 3'b111; end
            18'b100010011100111110: begin rgb_reg = 3'b111; end
            18'b100010011100111111: begin rgb_reg = 3'b111; end
            18'b100010011101000000: begin rgb_reg = 3'b111; end
            18'b100010011101000001: begin rgb_reg = 3'b111; end
            18'b100010011101000010: begin rgb_reg = 3'b111; end
            18'b100010100011000000: begin rgb_reg = 3'b111; end
            18'b100010100011000001: begin rgb_reg = 3'b111; end
            18'b100010100011000010: begin rgb_reg = 3'b111; end
            18'b100010100011000011: begin rgb_reg = 3'b111; end
            18'b100010100011000100: begin rgb_reg = 3'b111; end
            18'b100010100011000101: begin rgb_reg = 3'b111; end
            18'b100010100011000110: begin rgb_reg = 3'b111; end
            18'b100010100011001110: begin rgb_reg = 3'b111; end
            18'b100010100011001111: begin rgb_reg = 3'b111; end
            18'b100010100011010000: begin rgb_reg = 3'b111; end
            18'b100010100011010001: begin rgb_reg = 3'b111; end
            18'b100010100011010010: begin rgb_reg = 3'b111; end
            18'b100010100011010011: begin rgb_reg = 3'b111; end
            18'b100010100011011011: begin rgb_reg = 3'b111; end
            18'b100010100011011100: begin rgb_reg = 3'b111; end
            18'b100010100011011101: begin rgb_reg = 3'b111; end
            18'b100010100011011110: begin rgb_reg = 3'b111; end
            18'b100010100011011111: begin rgb_reg = 3'b111; end
            18'b100010100011100000: begin rgb_reg = 3'b111; end
            18'b100010100011100001: begin rgb_reg = 3'b111; end
            18'b100010100011101001: begin rgb_reg = 3'b111; end
            18'b100010100011101010: begin rgb_reg = 3'b111; end
            18'b100010100011101011: begin rgb_reg = 3'b111; end
            18'b100010100011101100: begin rgb_reg = 3'b111; end
            18'b100010100011101101: begin rgb_reg = 3'b111; end
            18'b100010100011101110: begin rgb_reg = 3'b111; end
            18'b100010100011110100: begin rgb_reg = 3'b111; end
            18'b100010100011110101: begin rgb_reg = 3'b111; end
            18'b100010100011110110: begin rgb_reg = 3'b111; end
            18'b100010100011110111: begin rgb_reg = 3'b111; end
            18'b100010100011111000: begin rgb_reg = 3'b111; end
            18'b100010100011111001: begin rgb_reg = 3'b111; end
            18'b100010100011111010: begin rgb_reg = 3'b111; end
            18'b100010100011111011: begin rgb_reg = 3'b111; end
            18'b100010100011111100: begin rgb_reg = 3'b111; end
            18'b100010100011111101: begin rgb_reg = 3'b111; end
            18'b100010100011111110: begin rgb_reg = 3'b111; end
            18'b100010100100000001: begin rgb_reg = 3'b111; end
            18'b100010100100000010: begin rgb_reg = 3'b111; end
            18'b100010100100000011: begin rgb_reg = 3'b111; end
            18'b100010100100000100: begin rgb_reg = 3'b111; end
            18'b100010100100000101: begin rgb_reg = 3'b111; end
            18'b100010100100000110: begin rgb_reg = 3'b111; end
            18'b100010100100000111: begin rgb_reg = 3'b111; end
            18'b100010100100001000: begin rgb_reg = 3'b111; end
            18'b100010100100001001: begin rgb_reg = 3'b111; end
            18'b100010100100001010: begin rgb_reg = 3'b111; end
            18'b100010100100001011: begin rgb_reg = 3'b111; end
            18'b100010100100010001: begin rgb_reg = 3'b111; end
            18'b100010100100010010: begin rgb_reg = 3'b111; end
            18'b100010100100010011: begin rgb_reg = 3'b111; end
            18'b100010100100010100: begin rgb_reg = 3'b111; end
            18'b100010100100010101: begin rgb_reg = 3'b111; end
            18'b100010100100010110: begin rgb_reg = 3'b111; end
            18'b100010100100010111: begin rgb_reg = 3'b111; end
            18'b100010100100011100: begin rgb_reg = 3'b111; end
            18'b100010100100011101: begin rgb_reg = 3'b111; end
            18'b100010100100011110: begin rgb_reg = 3'b111; end
            18'b100010100100011111: begin rgb_reg = 3'b111; end
            18'b100010100100100000: begin rgb_reg = 3'b111; end
            18'b100010100100100001: begin rgb_reg = 3'b111; end
            18'b100010100100100010: begin rgb_reg = 3'b111; end
            18'b100010100100100011: begin rgb_reg = 3'b111; end
            18'b100010100100100100: begin rgb_reg = 3'b111; end
            18'b100010100100100101: begin rgb_reg = 3'b111; end
            18'b100010100100100110: begin rgb_reg = 3'b111; end
            18'b100010100100101010: begin rgb_reg = 3'b111; end
            18'b100010100100101011: begin rgb_reg = 3'b111; end
            18'b100010100100101100: begin rgb_reg = 3'b111; end
            18'b100010100100101101: begin rgb_reg = 3'b111; end
            18'b100010100100101110: begin rgb_reg = 3'b111; end
            18'b100010100100101111: begin rgb_reg = 3'b111; end
            18'b100010100100110000: begin rgb_reg = 3'b111; end
            18'b100010100100110001: begin rgb_reg = 3'b111; end
            18'b100010100100110010: begin rgb_reg = 3'b111; end
            18'b100010100100110011: begin rgb_reg = 3'b111; end
            18'b100010100100110100: begin rgb_reg = 3'b111; end
            18'b100010100100110111: begin rgb_reg = 3'b111; end
            18'b100010100100111000: begin rgb_reg = 3'b111; end
            18'b100010100100111001: begin rgb_reg = 3'b111; end
            18'b100010100100111010: begin rgb_reg = 3'b111; end
            18'b100010100100111011: begin rgb_reg = 3'b111; end
            18'b100010100100111100: begin rgb_reg = 3'b111; end
            18'b100010100100111101: begin rgb_reg = 3'b111; end
            18'b100010100100111110: begin rgb_reg = 3'b111; end
            18'b100010100100111111: begin rgb_reg = 3'b111; end
            18'b100010100101000000: begin rgb_reg = 3'b111; end
            18'b100010100101000001: begin rgb_reg = 3'b111; end
            18'b100011011001110111: begin rgb_reg = 3'b111; end
            18'b100011011001111000: begin rgb_reg = 3'b111; end
            18'b100011011001111001: begin rgb_reg = 3'b111; end
            18'b100011011001111010: begin rgb_reg = 3'b111; end
            18'b100011011001111011: begin rgb_reg = 3'b111; end
            18'b100011011001111100: begin rgb_reg = 3'b111; end
            18'b100011011001111101: begin rgb_reg = 3'b111; end
            18'b100011011001111110: begin rgb_reg = 3'b111; end
            18'b100011011001111111: begin rgb_reg = 3'b111; end
            18'b100011011010000000: begin rgb_reg = 3'b111; end
            18'b100011011010000011: begin rgb_reg = 3'b111; end
            18'b100011011010000100: begin rgb_reg = 3'b111; end
            18'b100011011011010111: begin rgb_reg = 3'b111; end
            18'b100011011011011000: begin rgb_reg = 3'b111; end
            18'b100011011011011111: begin rgb_reg = 3'b111; end
            18'b100011011011100000: begin rgb_reg = 3'b111; end
            18'b100011011100110111: begin rgb_reg = 3'b111; end
            18'b100011011100111000: begin rgb_reg = 3'b111; end
            18'b100011011101010011: begin rgb_reg = 3'b111; end
            18'b100011011101010100: begin rgb_reg = 3'b111; end
            18'b100011011110000101: begin rgb_reg = 3'b111; end
            18'b100011011110000110: begin rgb_reg = 3'b111; end
            18'b100011100001110111: begin rgb_reg = 3'b111; end
            18'b100011100001111000: begin rgb_reg = 3'b111; end
            18'b100011100001111001: begin rgb_reg = 3'b111; end
            18'b100011100001111010: begin rgb_reg = 3'b111; end
            18'b100011100001111011: begin rgb_reg = 3'b111; end
            18'b100011100001111100: begin rgb_reg = 3'b111; end
            18'b100011100001111101: begin rgb_reg = 3'b111; end
            18'b100011100001111110: begin rgb_reg = 3'b111; end
            18'b100011100001111111: begin rgb_reg = 3'b111; end
            18'b100011100010000000: begin rgb_reg = 3'b111; end
            18'b100011100010000011: begin rgb_reg = 3'b111; end
            18'b100011100010000100: begin rgb_reg = 3'b111; end
            18'b100011100011010111: begin rgb_reg = 3'b111; end
            18'b100011100011011000: begin rgb_reg = 3'b111; end
            18'b100011100011011111: begin rgb_reg = 3'b111; end
            18'b100011100011100000: begin rgb_reg = 3'b111; end
            18'b100011100100110111: begin rgb_reg = 3'b111; end
            18'b100011100100111000: begin rgb_reg = 3'b111; end
            18'b100011100101010011: begin rgb_reg = 3'b111; end
            18'b100011100101010100: begin rgb_reg = 3'b111; end
            18'b100011100110000101: begin rgb_reg = 3'b111; end
            18'b100011100110000110: begin rgb_reg = 3'b111; end
            18'b100011101001111011: begin rgb_reg = 3'b111; end
            18'b100011101001111100: begin rgb_reg = 3'b111; end
            18'b100011101010000011: begin rgb_reg = 3'b111; end
            18'b100011101010000100: begin rgb_reg = 3'b111; end
            18'b100011101011010111: begin rgb_reg = 3'b111; end
            18'b100011101011011000: begin rgb_reg = 3'b111; end
            18'b100011101011011101: begin rgb_reg = 3'b111; end
            18'b100011101011011110: begin rgb_reg = 3'b111; end
            18'b100011101101010011: begin rgb_reg = 3'b111; end
            18'b100011101101010100: begin rgb_reg = 3'b111; end
            18'b100011101110000011: begin rgb_reg = 3'b111; end
            18'b100011101110000100: begin rgb_reg = 3'b111; end
            18'b100011101110000101: begin rgb_reg = 3'b111; end
            18'b100011101110000110: begin rgb_reg = 3'b111; end
            18'b100011101110000111: begin rgb_reg = 3'b111; end
            18'b100011101110001000: begin rgb_reg = 3'b111; end
            18'b100011110001111011: begin rgb_reg = 3'b111; end
            18'b100011110001111100: begin rgb_reg = 3'b111; end
            18'b100011110010000011: begin rgb_reg = 3'b111; end
            18'b100011110010000100: begin rgb_reg = 3'b111; end
            18'b100011110011010111: begin rgb_reg = 3'b111; end
            18'b100011110011011000: begin rgb_reg = 3'b111; end
            18'b100011110011011101: begin rgb_reg = 3'b111; end
            18'b100011110011011110: begin rgb_reg = 3'b111; end
            18'b100011110101010011: begin rgb_reg = 3'b111; end
            18'b100011110101010100: begin rgb_reg = 3'b111; end
            18'b100011110110000011: begin rgb_reg = 3'b111; end
            18'b100011110110000100: begin rgb_reg = 3'b111; end
            18'b100011110110000101: begin rgb_reg = 3'b111; end
            18'b100011110110000110: begin rgb_reg = 3'b111; end
            18'b100011110110000111: begin rgb_reg = 3'b111; end
            18'b100011110110001000: begin rgb_reg = 3'b111; end
            18'b100011111001111011: begin rgb_reg = 3'b111; end
            18'b100011111001111100: begin rgb_reg = 3'b111; end
            18'b100011111010000011: begin rgb_reg = 3'b111; end
            18'b100011111010000100: begin rgb_reg = 3'b111; end
            18'b100011111010000111: begin rgb_reg = 3'b111; end
            18'b100011111010001000: begin rgb_reg = 3'b111; end
            18'b100011111010001001: begin rgb_reg = 3'b111; end
            18'b100011111010001010: begin rgb_reg = 3'b111; end
            18'b100011111010010001: begin rgb_reg = 3'b111; end
            18'b100011111010010010: begin rgb_reg = 3'b111; end
            18'b100011111010010011: begin rgb_reg = 3'b111; end
            18'b100011111010010100: begin rgb_reg = 3'b111; end
            18'b100011111010010101: begin rgb_reg = 3'b111; end
            18'b100011111010010110: begin rgb_reg = 3'b111; end
            18'b100011111010011011: begin rgb_reg = 3'b111; end
            18'b100011111010011100: begin rgb_reg = 3'b111; end
            18'b100011111010100011: begin rgb_reg = 3'b111; end
            18'b100011111010100100: begin rgb_reg = 3'b111; end
            18'b100011111010101001: begin rgb_reg = 3'b111; end
            18'b100011111010101010: begin rgb_reg = 3'b111; end
            18'b100011111010101011: begin rgb_reg = 3'b111; end
            18'b100011111010101100: begin rgb_reg = 3'b111; end
            18'b100011111010101101: begin rgb_reg = 3'b111; end
            18'b100011111010101110: begin rgb_reg = 3'b111; end
            18'b100011111010110011: begin rgb_reg = 3'b111; end
            18'b100011111010110100: begin rgb_reg = 3'b111; end
            18'b100011111010110111: begin rgb_reg = 3'b111; end
            18'b100011111010111000: begin rgb_reg = 3'b111; end
            18'b100011111010111001: begin rgb_reg = 3'b111; end
            18'b100011111010111010: begin rgb_reg = 3'b111; end
            18'b100011111010111111: begin rgb_reg = 3'b111; end
            18'b100011111011000000: begin rgb_reg = 3'b111; end
            18'b100011111011000001: begin rgb_reg = 3'b111; end
            18'b100011111011000010: begin rgb_reg = 3'b111; end
            18'b100011111011000011: begin rgb_reg = 3'b111; end
            18'b100011111011000100: begin rgb_reg = 3'b111; end
            18'b100011111011000101: begin rgb_reg = 3'b111; end
            18'b100011111011000110: begin rgb_reg = 3'b111; end
            18'b100011111011010111: begin rgb_reg = 3'b111; end
            18'b100011111011011000: begin rgb_reg = 3'b111; end
            18'b100011111011011001: begin rgb_reg = 3'b111; end
            18'b100011111011011010: begin rgb_reg = 3'b111; end
            18'b100011111011011011: begin rgb_reg = 3'b111; end
            18'b100011111011011100: begin rgb_reg = 3'b111; end
            18'b100011111011100101: begin rgb_reg = 3'b111; end
            18'b100011111011100110: begin rgb_reg = 3'b111; end
            18'b100011111011100111: begin rgb_reg = 3'b111; end
            18'b100011111011101000: begin rgb_reg = 3'b111; end
            18'b100011111011101001: begin rgb_reg = 3'b111; end
            18'b100011111011101010: begin rgb_reg = 3'b111; end
            18'b100011111011101111: begin rgb_reg = 3'b111; end
            18'b100011111011110000: begin rgb_reg = 3'b111; end
            18'b100011111011110001: begin rgb_reg = 3'b111; end
            18'b100011111011110010: begin rgb_reg = 3'b111; end
            18'b100011111011110011: begin rgb_reg = 3'b111; end
            18'b100011111011110100: begin rgb_reg = 3'b111; end
            18'b100011111011110101: begin rgb_reg = 3'b111; end
            18'b100011111011110110: begin rgb_reg = 3'b111; end
            18'b100011111011111101: begin rgb_reg = 3'b111; end
            18'b100011111011111110: begin rgb_reg = 3'b111; end
            18'b100011111011111111: begin rgb_reg = 3'b111; end
            18'b100011111100000000: begin rgb_reg = 3'b111; end
            18'b100011111100000001: begin rgb_reg = 3'b111; end
            18'b100011111100000010: begin rgb_reg = 3'b111; end
            18'b100011111100000011: begin rgb_reg = 3'b111; end
            18'b100011111100000100: begin rgb_reg = 3'b111; end
            18'b100011111100000111: begin rgb_reg = 3'b111; end
            18'b100011111100001000: begin rgb_reg = 3'b111; end
            18'b100011111100001111: begin rgb_reg = 3'b111; end
            18'b100011111100010000: begin rgb_reg = 3'b111; end
            18'b100011111100010101: begin rgb_reg = 3'b111; end
            18'b100011111100010110: begin rgb_reg = 3'b111; end
            18'b100011111100010111: begin rgb_reg = 3'b111; end
            18'b100011111100011000: begin rgb_reg = 3'b111; end
            18'b100011111100011001: begin rgb_reg = 3'b111; end
            18'b100011111100011010: begin rgb_reg = 3'b111; end
            18'b100011111100011111: begin rgb_reg = 3'b111; end
            18'b100011111100100000: begin rgb_reg = 3'b111; end
            18'b100011111100100001: begin rgb_reg = 3'b111; end
            18'b100011111100100010: begin rgb_reg = 3'b111; end
            18'b100011111100100011: begin rgb_reg = 3'b111; end
            18'b100011111100100100: begin rgb_reg = 3'b111; end
            18'b100011111100100101: begin rgb_reg = 3'b111; end
            18'b100011111100100110: begin rgb_reg = 3'b111; end
            18'b100011111100101101: begin rgb_reg = 3'b111; end
            18'b100011111100101110: begin rgb_reg = 3'b111; end
            18'b100011111100101111: begin rgb_reg = 3'b111; end
            18'b100011111100110000: begin rgb_reg = 3'b111; end
            18'b100011111100110001: begin rgb_reg = 3'b111; end
            18'b100011111100110010: begin rgb_reg = 3'b111; end
            18'b100011111100110011: begin rgb_reg = 3'b111; end
            18'b100011111100110100: begin rgb_reg = 3'b111; end
            18'b100011111100110111: begin rgb_reg = 3'b111; end
            18'b100011111100111000: begin rgb_reg = 3'b111; end
            18'b100011111100111011: begin rgb_reg = 3'b111; end
            18'b100011111100111100: begin rgb_reg = 3'b111; end
            18'b100011111100111101: begin rgb_reg = 3'b111; end
            18'b100011111100111110: begin rgb_reg = 3'b111; end
            18'b100011111100111111: begin rgb_reg = 3'b111; end
            18'b100011111101000000: begin rgb_reg = 3'b111; end
            18'b100011111101000001: begin rgb_reg = 3'b111; end
            18'b100011111101000010: begin rgb_reg = 3'b111; end
            18'b100011111101001001: begin rgb_reg = 3'b111; end
            18'b100011111101001010: begin rgb_reg = 3'b111; end
            18'b100011111101001011: begin rgb_reg = 3'b111; end
            18'b100011111101001100: begin rgb_reg = 3'b111; end
            18'b100011111101001101: begin rgb_reg = 3'b111; end
            18'b100011111101001110: begin rgb_reg = 3'b111; end
            18'b100011111101001111: begin rgb_reg = 3'b111; end
            18'b100011111101010000: begin rgb_reg = 3'b111; end
            18'b100011111101010011: begin rgb_reg = 3'b111; end
            18'b100011111101010100: begin rgb_reg = 3'b111; end
            18'b100011111101010111: begin rgb_reg = 3'b111; end
            18'b100011111101011000: begin rgb_reg = 3'b111; end
            18'b100011111101011001: begin rgb_reg = 3'b111; end
            18'b100011111101011010: begin rgb_reg = 3'b111; end
            18'b100011111101100001: begin rgb_reg = 3'b111; end
            18'b100011111101100010: begin rgb_reg = 3'b111; end
            18'b100011111101100011: begin rgb_reg = 3'b111; end
            18'b100011111101100100: begin rgb_reg = 3'b111; end
            18'b100011111101100101: begin rgb_reg = 3'b111; end
            18'b100011111101100110: begin rgb_reg = 3'b111; end
            18'b100011111101101011: begin rgb_reg = 3'b111; end
            18'b100011111101101100: begin rgb_reg = 3'b111; end
            18'b100011111101101101: begin rgb_reg = 3'b111; end
            18'b100011111101101110: begin rgb_reg = 3'b111; end
            18'b100011111101101111: begin rgb_reg = 3'b111; end
            18'b100011111101110000: begin rgb_reg = 3'b111; end
            18'b100011111101110001: begin rgb_reg = 3'b111; end
            18'b100011111101110010: begin rgb_reg = 3'b111; end
            18'b100011111101111001: begin rgb_reg = 3'b111; end
            18'b100011111101111010: begin rgb_reg = 3'b111; end
            18'b100011111101111011: begin rgb_reg = 3'b111; end
            18'b100011111101111100: begin rgb_reg = 3'b111; end
            18'b100011111101111101: begin rgb_reg = 3'b111; end
            18'b100011111101111110: begin rgb_reg = 3'b111; end
            18'b100011111110000101: begin rgb_reg = 3'b111; end
            18'b100011111110000110: begin rgb_reg = 3'b111; end
            18'b100100000001111011: begin rgb_reg = 3'b111; end
            18'b100100000001111100: begin rgb_reg = 3'b111; end
            18'b100100000010000011: begin rgb_reg = 3'b111; end
            18'b100100000010000100: begin rgb_reg = 3'b111; end
            18'b100100000010000111: begin rgb_reg = 3'b111; end
            18'b100100000010001000: begin rgb_reg = 3'b111; end
            18'b100100000010001001: begin rgb_reg = 3'b111; end
            18'b100100000010001010: begin rgb_reg = 3'b111; end
            18'b100100000010010001: begin rgb_reg = 3'b111; end
            18'b100100000010010010: begin rgb_reg = 3'b111; end
            18'b100100000010010011: begin rgb_reg = 3'b111; end
            18'b100100000010010100: begin rgb_reg = 3'b111; end
            18'b100100000010010101: begin rgb_reg = 3'b111; end
            18'b100100000010010110: begin rgb_reg = 3'b111; end
            18'b100100000010011011: begin rgb_reg = 3'b111; end
            18'b100100000010011100: begin rgb_reg = 3'b111; end
            18'b100100000010100011: begin rgb_reg = 3'b111; end
            18'b100100000010100100: begin rgb_reg = 3'b111; end
            18'b100100000010101001: begin rgb_reg = 3'b111; end
            18'b100100000010101010: begin rgb_reg = 3'b111; end
            18'b100100000010101011: begin rgb_reg = 3'b111; end
            18'b100100000010101100: begin rgb_reg = 3'b111; end
            18'b100100000010101101: begin rgb_reg = 3'b111; end
            18'b100100000010101110: begin rgb_reg = 3'b111; end
            18'b100100000010110011: begin rgb_reg = 3'b111; end
            18'b100100000010110100: begin rgb_reg = 3'b111; end
            18'b100100000010110111: begin rgb_reg = 3'b111; end
            18'b100100000010111000: begin rgb_reg = 3'b111; end
            18'b100100000010111001: begin rgb_reg = 3'b111; end
            18'b100100000010111010: begin rgb_reg = 3'b111; end
            18'b100100000010111111: begin rgb_reg = 3'b111; end
            18'b100100000011000000: begin rgb_reg = 3'b111; end
            18'b100100000011000001: begin rgb_reg = 3'b111; end
            18'b100100000011000010: begin rgb_reg = 3'b111; end
            18'b100100000011000011: begin rgb_reg = 3'b111; end
            18'b100100000011000100: begin rgb_reg = 3'b111; end
            18'b100100000011000101: begin rgb_reg = 3'b111; end
            18'b100100000011000110: begin rgb_reg = 3'b111; end
            18'b100100000011010111: begin rgb_reg = 3'b111; end
            18'b100100000011011000: begin rgb_reg = 3'b111; end
            18'b100100000011011001: begin rgb_reg = 3'b111; end
            18'b100100000011011010: begin rgb_reg = 3'b111; end
            18'b100100000011011011: begin rgb_reg = 3'b111; end
            18'b100100000011011100: begin rgb_reg = 3'b111; end
            18'b100100000011100101: begin rgb_reg = 3'b111; end
            18'b100100000011100110: begin rgb_reg = 3'b111; end
            18'b100100000011100111: begin rgb_reg = 3'b111; end
            18'b100100000011101000: begin rgb_reg = 3'b111; end
            18'b100100000011101001: begin rgb_reg = 3'b111; end
            18'b100100000011101010: begin rgb_reg = 3'b111; end
            18'b100100000011101111: begin rgb_reg = 3'b111; end
            18'b100100000011110000: begin rgb_reg = 3'b111; end
            18'b100100000011110001: begin rgb_reg = 3'b111; end
            18'b100100000011110010: begin rgb_reg = 3'b111; end
            18'b100100000011110011: begin rgb_reg = 3'b111; end
            18'b100100000011110100: begin rgb_reg = 3'b111; end
            18'b100100000011110101: begin rgb_reg = 3'b111; end
            18'b100100000011110110: begin rgb_reg = 3'b111; end
            18'b100100000011111101: begin rgb_reg = 3'b111; end
            18'b100100000011111110: begin rgb_reg = 3'b111; end
            18'b100100000011111111: begin rgb_reg = 3'b111; end
            18'b100100000100000000: begin rgb_reg = 3'b111; end
            18'b100100000100000001: begin rgb_reg = 3'b111; end
            18'b100100000100000010: begin rgb_reg = 3'b111; end
            18'b100100000100000011: begin rgb_reg = 3'b111; end
            18'b100100000100000100: begin rgb_reg = 3'b111; end
            18'b100100000100000111: begin rgb_reg = 3'b111; end
            18'b100100000100001000: begin rgb_reg = 3'b111; end
            18'b100100000100001111: begin rgb_reg = 3'b111; end
            18'b100100000100010000: begin rgb_reg = 3'b111; end
            18'b100100000100010101: begin rgb_reg = 3'b111; end
            18'b100100000100010110: begin rgb_reg = 3'b111; end
            18'b100100000100010111: begin rgb_reg = 3'b111; end
            18'b100100000100011000: begin rgb_reg = 3'b111; end
            18'b100100000100011001: begin rgb_reg = 3'b111; end
            18'b100100000100011010: begin rgb_reg = 3'b111; end
            18'b100100000100011111: begin rgb_reg = 3'b111; end
            18'b100100000100100000: begin rgb_reg = 3'b111; end
            18'b100100000100100001: begin rgb_reg = 3'b111; end
            18'b100100000100100010: begin rgb_reg = 3'b111; end
            18'b100100000100100011: begin rgb_reg = 3'b111; end
            18'b100100000100100100: begin rgb_reg = 3'b111; end
            18'b100100000100100101: begin rgb_reg = 3'b111; end
            18'b100100000100100110: begin rgb_reg = 3'b111; end
            18'b100100000100101101: begin rgb_reg = 3'b111; end
            18'b100100000100101110: begin rgb_reg = 3'b111; end
            18'b100100000100101111: begin rgb_reg = 3'b111; end
            18'b100100000100110000: begin rgb_reg = 3'b111; end
            18'b100100000100110001: begin rgb_reg = 3'b111; end
            18'b100100000100110010: begin rgb_reg = 3'b111; end
            18'b100100000100110011: begin rgb_reg = 3'b111; end
            18'b100100000100110100: begin rgb_reg = 3'b111; end
            18'b100100000100110111: begin rgb_reg = 3'b111; end
            18'b100100000100111000: begin rgb_reg = 3'b111; end
            18'b100100000100111011: begin rgb_reg = 3'b111; end
            18'b100100000100111100: begin rgb_reg = 3'b111; end
            18'b100100000100111101: begin rgb_reg = 3'b111; end
            18'b100100000100111110: begin rgb_reg = 3'b111; end
            18'b100100000100111111: begin rgb_reg = 3'b111; end
            18'b100100000101000000: begin rgb_reg = 3'b111; end
            18'b100100000101000001: begin rgb_reg = 3'b111; end
            18'b100100000101000010: begin rgb_reg = 3'b111; end
            18'b100100000101001001: begin rgb_reg = 3'b111; end
            18'b100100000101001010: begin rgb_reg = 3'b111; end
            18'b100100000101001011: begin rgb_reg = 3'b111; end
            18'b100100000101001100: begin rgb_reg = 3'b111; end
            18'b100100000101001101: begin rgb_reg = 3'b111; end
            18'b100100000101001110: begin rgb_reg = 3'b111; end
            18'b100100000101001111: begin rgb_reg = 3'b111; end
            18'b100100000101010000: begin rgb_reg = 3'b111; end
            18'b100100000101010011: begin rgb_reg = 3'b111; end
            18'b100100000101010100: begin rgb_reg = 3'b111; end
            18'b100100000101010111: begin rgb_reg = 3'b111; end
            18'b100100000101011000: begin rgb_reg = 3'b111; end
            18'b100100000101011001: begin rgb_reg = 3'b111; end
            18'b100100000101011010: begin rgb_reg = 3'b111; end
            18'b100100000101100001: begin rgb_reg = 3'b111; end
            18'b100100000101100010: begin rgb_reg = 3'b111; end
            18'b100100000101100011: begin rgb_reg = 3'b111; end
            18'b100100000101100100: begin rgb_reg = 3'b111; end
            18'b100100000101100101: begin rgb_reg = 3'b111; end
            18'b100100000101100110: begin rgb_reg = 3'b111; end
            18'b100100000101101011: begin rgb_reg = 3'b111; end
            18'b100100000101101100: begin rgb_reg = 3'b111; end
            18'b100100000101101101: begin rgb_reg = 3'b111; end
            18'b100100000101101110: begin rgb_reg = 3'b111; end
            18'b100100000101101111: begin rgb_reg = 3'b111; end
            18'b100100000101110000: begin rgb_reg = 3'b111; end
            18'b100100000101110001: begin rgb_reg = 3'b111; end
            18'b100100000101110010: begin rgb_reg = 3'b111; end
            18'b100100000101111001: begin rgb_reg = 3'b111; end
            18'b100100000101111010: begin rgb_reg = 3'b111; end
            18'b100100000101111011: begin rgb_reg = 3'b111; end
            18'b100100000101111100: begin rgb_reg = 3'b111; end
            18'b100100000101111101: begin rgb_reg = 3'b111; end
            18'b100100000101111110: begin rgb_reg = 3'b111; end
            18'b100100000110000101: begin rgb_reg = 3'b111; end
            18'b100100000110000110: begin rgb_reg = 3'b111; end
            18'b100100001001111011: begin rgb_reg = 3'b111; end
            18'b100100001001111100: begin rgb_reg = 3'b111; end
            18'b100100001010000011: begin rgb_reg = 3'b111; end
            18'b100100001010000100: begin rgb_reg = 3'b111; end
            18'b100100001010000101: begin rgb_reg = 3'b111; end
            18'b100100001010000110: begin rgb_reg = 3'b111; end
            18'b100100001010001011: begin rgb_reg = 3'b111; end
            18'b100100001010001100: begin rgb_reg = 3'b111; end
            18'b100100001010010111: begin rgb_reg = 3'b111; end
            18'b100100001010011000: begin rgb_reg = 3'b111; end
            18'b100100001010011011: begin rgb_reg = 3'b111; end
            18'b100100001010011100: begin rgb_reg = 3'b111; end
            18'b100100001010100011: begin rgb_reg = 3'b111; end
            18'b100100001010100100: begin rgb_reg = 3'b111; end
            18'b100100001010100111: begin rgb_reg = 3'b111; end
            18'b100100001010101000: begin rgb_reg = 3'b111; end
            18'b100100001010101111: begin rgb_reg = 3'b111; end
            18'b100100001010110000: begin rgb_reg = 3'b111; end
            18'b100100001010110011: begin rgb_reg = 3'b111; end
            18'b100100001010110100: begin rgb_reg = 3'b111; end
            18'b100100001010110101: begin rgb_reg = 3'b111; end
            18'b100100001010110110: begin rgb_reg = 3'b111; end
            18'b100100001010111011: begin rgb_reg = 3'b111; end
            18'b100100001010111100: begin rgb_reg = 3'b111; end
            18'b100100001010111111: begin rgb_reg = 3'b111; end
            18'b100100001011000000: begin rgb_reg = 3'b111; end
            18'b100100001011000111: begin rgb_reg = 3'b111; end
            18'b100100001011001000: begin rgb_reg = 3'b111; end
            18'b100100001011010111: begin rgb_reg = 3'b111; end
            18'b100100001011011000: begin rgb_reg = 3'b111; end
            18'b100100001011011101: begin rgb_reg = 3'b111; end
            18'b100100001011011110: begin rgb_reg = 3'b111; end
            18'b100100001011101011: begin rgb_reg = 3'b111; end
            18'b100100001011101100: begin rgb_reg = 3'b111; end
            18'b100100001011101111: begin rgb_reg = 3'b111; end
            18'b100100001011110000: begin rgb_reg = 3'b111; end
            18'b100100001011110111: begin rgb_reg = 3'b111; end
            18'b100100001011111000: begin rgb_reg = 3'b111; end
            18'b100100001011111011: begin rgb_reg = 3'b111; end
            18'b100100001011111100: begin rgb_reg = 3'b111; end
            18'b100100001100000011: begin rgb_reg = 3'b111; end
            18'b100100001100000100: begin rgb_reg = 3'b111; end
            18'b100100001100000111: begin rgb_reg = 3'b111; end
            18'b100100001100001000: begin rgb_reg = 3'b111; end
            18'b100100001100001111: begin rgb_reg = 3'b111; end
            18'b100100001100010000: begin rgb_reg = 3'b111; end
            18'b100100001100011011: begin rgb_reg = 3'b111; end
            18'b100100001100011100: begin rgb_reg = 3'b111; end
            18'b100100001100011111: begin rgb_reg = 3'b111; end
            18'b100100001100100000: begin rgb_reg = 3'b111; end
            18'b100100001100100111: begin rgb_reg = 3'b111; end
            18'b100100001100101000: begin rgb_reg = 3'b111; end
            18'b100100001100101011: begin rgb_reg = 3'b111; end
            18'b100100001100101100: begin rgb_reg = 3'b111; end
            18'b100100001100110111: begin rgb_reg = 3'b111; end
            18'b100100001100111000: begin rgb_reg = 3'b111; end
            18'b100100001100111011: begin rgb_reg = 3'b111; end
            18'b100100001100111100: begin rgb_reg = 3'b111; end
            18'b100100001101000011: begin rgb_reg = 3'b111; end
            18'b100100001101000100: begin rgb_reg = 3'b111; end
            18'b100100001101000111: begin rgb_reg = 3'b111; end
            18'b100100001101001000: begin rgb_reg = 3'b111; end
            18'b100100001101001111: begin rgb_reg = 3'b111; end
            18'b100100001101010000: begin rgb_reg = 3'b111; end
            18'b100100001101010011: begin rgb_reg = 3'b111; end
            18'b100100001101010100: begin rgb_reg = 3'b111; end
            18'b100100001101010101: begin rgb_reg = 3'b111; end
            18'b100100001101010110: begin rgb_reg = 3'b111; end
            18'b100100001101011011: begin rgb_reg = 3'b111; end
            18'b100100001101011100: begin rgb_reg = 3'b111; end
            18'b100100001101100111: begin rgb_reg = 3'b111; end
            18'b100100001101101000: begin rgb_reg = 3'b111; end
            18'b100100001101101011: begin rgb_reg = 3'b111; end
            18'b100100001101101100: begin rgb_reg = 3'b111; end
            18'b100100001101110011: begin rgb_reg = 3'b111; end
            18'b100100001101110100: begin rgb_reg = 3'b111; end
            18'b100100001101111111: begin rgb_reg = 3'b111; end
            18'b100100001110000000: begin rgb_reg = 3'b111; end
            18'b100100001110000101: begin rgb_reg = 3'b111; end
            18'b100100001110000110: begin rgb_reg = 3'b111; end
            18'b100100010001111011: begin rgb_reg = 3'b111; end
            18'b100100010001111100: begin rgb_reg = 3'b111; end
            18'b100100010010000011: begin rgb_reg = 3'b111; end
            18'b100100010010000100: begin rgb_reg = 3'b111; end
            18'b100100010010000101: begin rgb_reg = 3'b111; end
            18'b100100010010000110: begin rgb_reg = 3'b111; end
            18'b100100010010001011: begin rgb_reg = 3'b111; end
            18'b100100010010001100: begin rgb_reg = 3'b111; end
            18'b100100010010010111: begin rgb_reg = 3'b111; end
            18'b100100010010011000: begin rgb_reg = 3'b111; end
            18'b100100010010011011: begin rgb_reg = 3'b111; end
            18'b100100010010011100: begin rgb_reg = 3'b111; end
            18'b100100010010100011: begin rgb_reg = 3'b111; end
            18'b100100010010100100: begin rgb_reg = 3'b111; end
            18'b100100010010100111: begin rgb_reg = 3'b111; end
            18'b100100010010101000: begin rgb_reg = 3'b111; end
            18'b100100010010101111: begin rgb_reg = 3'b111; end
            18'b100100010010110000: begin rgb_reg = 3'b111; end
            18'b100100010010110011: begin rgb_reg = 3'b111; end
            18'b100100010010110100: begin rgb_reg = 3'b111; end
            18'b100100010010110101: begin rgb_reg = 3'b111; end
            18'b100100010010110110: begin rgb_reg = 3'b111; end
            18'b100100010010111011: begin rgb_reg = 3'b111; end
            18'b100100010010111100: begin rgb_reg = 3'b111; end
            18'b100100010010111111: begin rgb_reg = 3'b111; end
            18'b100100010011000000: begin rgb_reg = 3'b111; end
            18'b100100010011000111: begin rgb_reg = 3'b111; end
            18'b100100010011001000: begin rgb_reg = 3'b111; end
            18'b100100010011010111: begin rgb_reg = 3'b111; end
            18'b100100010011011000: begin rgb_reg = 3'b111; end
            18'b100100010011011101: begin rgb_reg = 3'b111; end
            18'b100100010011011110: begin rgb_reg = 3'b111; end
            18'b100100010011101011: begin rgb_reg = 3'b111; end
            18'b100100010011101100: begin rgb_reg = 3'b111; end
            18'b100100010011101111: begin rgb_reg = 3'b111; end
            18'b100100010011110000: begin rgb_reg = 3'b111; end
            18'b100100010011110111: begin rgb_reg = 3'b111; end
            18'b100100010011111000: begin rgb_reg = 3'b111; end
            18'b100100010011111011: begin rgb_reg = 3'b111; end
            18'b100100010011111100: begin rgb_reg = 3'b111; end
            18'b100100010100000011: begin rgb_reg = 3'b111; end
            18'b100100010100000100: begin rgb_reg = 3'b111; end
            18'b100100010100000111: begin rgb_reg = 3'b111; end
            18'b100100010100001000: begin rgb_reg = 3'b111; end
            18'b100100010100001111: begin rgb_reg = 3'b111; end
            18'b100100010100010000: begin rgb_reg = 3'b111; end
            18'b100100010100011011: begin rgb_reg = 3'b111; end
            18'b100100010100011100: begin rgb_reg = 3'b111; end
            18'b100100010100011111: begin rgb_reg = 3'b111; end
            18'b100100010100100000: begin rgb_reg = 3'b111; end
            18'b100100010100100111: begin rgb_reg = 3'b111; end
            18'b100100010100101000: begin rgb_reg = 3'b111; end
            18'b100100010100101011: begin rgb_reg = 3'b111; end
            18'b100100010100101100: begin rgb_reg = 3'b111; end
            18'b100100010100110111: begin rgb_reg = 3'b111; end
            18'b100100010100111000: begin rgb_reg = 3'b111; end
            18'b100100010100111011: begin rgb_reg = 3'b111; end
            18'b100100010100111100: begin rgb_reg = 3'b111; end
            18'b100100010101000011: begin rgb_reg = 3'b111; end
            18'b100100010101000100: begin rgb_reg = 3'b111; end
            18'b100100010101000111: begin rgb_reg = 3'b111; end
            18'b100100010101001000: begin rgb_reg = 3'b111; end
            18'b100100010101001111: begin rgb_reg = 3'b111; end
            18'b100100010101010000: begin rgb_reg = 3'b111; end
            18'b100100010101010011: begin rgb_reg = 3'b111; end
            18'b100100010101010100: begin rgb_reg = 3'b111; end
            18'b100100010101010101: begin rgb_reg = 3'b111; end
            18'b100100010101010110: begin rgb_reg = 3'b111; end
            18'b100100010101011011: begin rgb_reg = 3'b111; end
            18'b100100010101011100: begin rgb_reg = 3'b111; end
            18'b100100010101100111: begin rgb_reg = 3'b111; end
            18'b100100010101101000: begin rgb_reg = 3'b111; end
            18'b100100010101101011: begin rgb_reg = 3'b111; end
            18'b100100010101101100: begin rgb_reg = 3'b111; end
            18'b100100010101110011: begin rgb_reg = 3'b111; end
            18'b100100010101110100: begin rgb_reg = 3'b111; end
            18'b100100010101111111: begin rgb_reg = 3'b111; end
            18'b100100010110000000: begin rgb_reg = 3'b111; end
            18'b100100010110000101: begin rgb_reg = 3'b111; end
            18'b100100010110000110: begin rgb_reg = 3'b111; end
            18'b100100011001111011: begin rgb_reg = 3'b111; end
            18'b100100011001111100: begin rgb_reg = 3'b111; end
            18'b100100011010000011: begin rgb_reg = 3'b111; end
            18'b100100011010000100: begin rgb_reg = 3'b111; end
            18'b100100011010001011: begin rgb_reg = 3'b111; end
            18'b100100011010001100: begin rgb_reg = 3'b111; end
            18'b100100011010010001: begin rgb_reg = 3'b111; end
            18'b100100011010010010: begin rgb_reg = 3'b111; end
            18'b100100011010010011: begin rgb_reg = 3'b111; end
            18'b100100011010010100: begin rgb_reg = 3'b111; end
            18'b100100011010010101: begin rgb_reg = 3'b111; end
            18'b100100011010010110: begin rgb_reg = 3'b111; end
            18'b100100011010010111: begin rgb_reg = 3'b111; end
            18'b100100011010011000: begin rgb_reg = 3'b111; end
            18'b100100011010011011: begin rgb_reg = 3'b111; end
            18'b100100011010011100: begin rgb_reg = 3'b111; end
            18'b100100011010011111: begin rgb_reg = 3'b111; end
            18'b100100011010100000: begin rgb_reg = 3'b111; end
            18'b100100011010100011: begin rgb_reg = 3'b111; end
            18'b100100011010100100: begin rgb_reg = 3'b111; end
            18'b100100011010100111: begin rgb_reg = 3'b111; end
            18'b100100011010101000: begin rgb_reg = 3'b111; end
            18'b100100011010101111: begin rgb_reg = 3'b111; end
            18'b100100011010110000: begin rgb_reg = 3'b111; end
            18'b100100011010110011: begin rgb_reg = 3'b111; end
            18'b100100011010110100: begin rgb_reg = 3'b111; end
            18'b100100011010111111: begin rgb_reg = 3'b111; end
            18'b100100011011000000: begin rgb_reg = 3'b111; end
            18'b100100011011000111: begin rgb_reg = 3'b111; end
            18'b100100011011001000: begin rgb_reg = 3'b111; end
            18'b100100011011010111: begin rgb_reg = 3'b111; end
            18'b100100011011011000: begin rgb_reg = 3'b111; end
            18'b100100011011011111: begin rgb_reg = 3'b111; end
            18'b100100011011100000: begin rgb_reg = 3'b111; end
            18'b100100011011100101: begin rgb_reg = 3'b111; end
            18'b100100011011100110: begin rgb_reg = 3'b111; end
            18'b100100011011100111: begin rgb_reg = 3'b111; end
            18'b100100011011101000: begin rgb_reg = 3'b111; end
            18'b100100011011101001: begin rgb_reg = 3'b111; end
            18'b100100011011101010: begin rgb_reg = 3'b111; end
            18'b100100011011101011: begin rgb_reg = 3'b111; end
            18'b100100011011101100: begin rgb_reg = 3'b111; end
            18'b100100011011101111: begin rgb_reg = 3'b111; end
            18'b100100011011110000: begin rgb_reg = 3'b111; end
            18'b100100011011110111: begin rgb_reg = 3'b111; end
            18'b100100011011111000: begin rgb_reg = 3'b111; end
            18'b100100011011111011: begin rgb_reg = 3'b111; end
            18'b100100011011111100: begin rgb_reg = 3'b111; end
            18'b100100011100000011: begin rgb_reg = 3'b111; end
            18'b100100011100000100: begin rgb_reg = 3'b111; end
            18'b100100011100000111: begin rgb_reg = 3'b111; end
            18'b100100011100001000: begin rgb_reg = 3'b111; end
            18'b100100011100001011: begin rgb_reg = 3'b111; end
            18'b100100011100001100: begin rgb_reg = 3'b111; end
            18'b100100011100001111: begin rgb_reg = 3'b111; end
            18'b100100011100010000: begin rgb_reg = 3'b111; end
            18'b100100011100010101: begin rgb_reg = 3'b111; end
            18'b100100011100010110: begin rgb_reg = 3'b111; end
            18'b100100011100010111: begin rgb_reg = 3'b111; end
            18'b100100011100011000: begin rgb_reg = 3'b111; end
            18'b100100011100011001: begin rgb_reg = 3'b111; end
            18'b100100011100011010: begin rgb_reg = 3'b111; end
            18'b100100011100011011: begin rgb_reg = 3'b111; end
            18'b100100011100011100: begin rgb_reg = 3'b111; end
            18'b100100011100011111: begin rgb_reg = 3'b111; end
            18'b100100011100100000: begin rgb_reg = 3'b111; end
            18'b100100011100100111: begin rgb_reg = 3'b111; end
            18'b100100011100101000: begin rgb_reg = 3'b111; end
            18'b100100011100101101: begin rgb_reg = 3'b111; end
            18'b100100011100101110: begin rgb_reg = 3'b111; end
            18'b100100011100101111: begin rgb_reg = 3'b111; end
            18'b100100011100110000: begin rgb_reg = 3'b111; end
            18'b100100011100110001: begin rgb_reg = 3'b111; end
            18'b100100011100110010: begin rgb_reg = 3'b111; end
            18'b100100011100110111: begin rgb_reg = 3'b111; end
            18'b100100011100111000: begin rgb_reg = 3'b111; end
            18'b100100011100111011: begin rgb_reg = 3'b111; end
            18'b100100011100111100: begin rgb_reg = 3'b111; end
            18'b100100011101000011: begin rgb_reg = 3'b111; end
            18'b100100011101000100: begin rgb_reg = 3'b111; end
            18'b100100011101000111: begin rgb_reg = 3'b111; end
            18'b100100011101001000: begin rgb_reg = 3'b111; end
            18'b100100011101001111: begin rgb_reg = 3'b111; end
            18'b100100011101010000: begin rgb_reg = 3'b111; end
            18'b100100011101010011: begin rgb_reg = 3'b111; end
            18'b100100011101010100: begin rgb_reg = 3'b111; end
            18'b100100011101011011: begin rgb_reg = 3'b111; end
            18'b100100011101011100: begin rgb_reg = 3'b111; end
            18'b100100011101100001: begin rgb_reg = 3'b111; end
            18'b100100011101100010: begin rgb_reg = 3'b111; end
            18'b100100011101100011: begin rgb_reg = 3'b111; end
            18'b100100011101100100: begin rgb_reg = 3'b111; end
            18'b100100011101100101: begin rgb_reg = 3'b111; end
            18'b100100011101100110: begin rgb_reg = 3'b111; end
            18'b100100011101100111: begin rgb_reg = 3'b111; end
            18'b100100011101101000: begin rgb_reg = 3'b111; end
            18'b100100011101101011: begin rgb_reg = 3'b111; end
            18'b100100011101101100: begin rgb_reg = 3'b111; end
            18'b100100011101110011: begin rgb_reg = 3'b111; end
            18'b100100011101110100: begin rgb_reg = 3'b111; end
            18'b100100011101111001: begin rgb_reg = 3'b111; end
            18'b100100011101111010: begin rgb_reg = 3'b111; end
            18'b100100011101111011: begin rgb_reg = 3'b111; end
            18'b100100011101111100: begin rgb_reg = 3'b111; end
            18'b100100011101111101: begin rgb_reg = 3'b111; end
            18'b100100011101111110: begin rgb_reg = 3'b111; end
            18'b100100011101111111: begin rgb_reg = 3'b111; end
            18'b100100011110000000: begin rgb_reg = 3'b111; end
            18'b100100011110000101: begin rgb_reg = 3'b111; end
            18'b100100011110000110: begin rgb_reg = 3'b111; end
            18'b100100100001111011: begin rgb_reg = 3'b111; end
            18'b100100100001111100: begin rgb_reg = 3'b111; end
            18'b100100100010000011: begin rgb_reg = 3'b111; end
            18'b100100100010000100: begin rgb_reg = 3'b111; end
            18'b100100100010001011: begin rgb_reg = 3'b111; end
            18'b100100100010001100: begin rgb_reg = 3'b111; end
            18'b100100100010010001: begin rgb_reg = 3'b111; end
            18'b100100100010010010: begin rgb_reg = 3'b111; end
            18'b100100100010010011: begin rgb_reg = 3'b111; end
            18'b100100100010010100: begin rgb_reg = 3'b111; end
            18'b100100100010010101: begin rgb_reg = 3'b111; end
            18'b100100100010010110: begin rgb_reg = 3'b111; end
            18'b100100100010010111: begin rgb_reg = 3'b111; end
            18'b100100100010011000: begin rgb_reg = 3'b111; end
            18'b100100100010011011: begin rgb_reg = 3'b111; end
            18'b100100100010011100: begin rgb_reg = 3'b111; end
            18'b100100100010011111: begin rgb_reg = 3'b111; end
            18'b100100100010100000: begin rgb_reg = 3'b111; end
            18'b100100100010100011: begin rgb_reg = 3'b111; end
            18'b100100100010100100: begin rgb_reg = 3'b111; end
            18'b100100100010100111: begin rgb_reg = 3'b111; end
            18'b100100100010101000: begin rgb_reg = 3'b111; end
            18'b100100100010101111: begin rgb_reg = 3'b111; end
            18'b100100100010110000: begin rgb_reg = 3'b111; end
            18'b100100100010110011: begin rgb_reg = 3'b111; end
            18'b100100100010110100: begin rgb_reg = 3'b111; end
            18'b100100100010111111: begin rgb_reg = 3'b111; end
            18'b100100100011000000: begin rgb_reg = 3'b111; end
            18'b100100100011000111: begin rgb_reg = 3'b111; end
            18'b100100100011001000: begin rgb_reg = 3'b111; end
            18'b100100100011010111: begin rgb_reg = 3'b111; end
            18'b100100100011011000: begin rgb_reg = 3'b111; end
            18'b100100100011011111: begin rgb_reg = 3'b111; end
            18'b100100100011100000: begin rgb_reg = 3'b111; end
            18'b100100100011100101: begin rgb_reg = 3'b111; end
            18'b100100100011100110: begin rgb_reg = 3'b111; end
            18'b100100100011100111: begin rgb_reg = 3'b111; end
            18'b100100100011101000: begin rgb_reg = 3'b111; end
            18'b100100100011101001: begin rgb_reg = 3'b111; end
            18'b100100100011101010: begin rgb_reg = 3'b111; end
            18'b100100100011101011: begin rgb_reg = 3'b111; end
            18'b100100100011101100: begin rgb_reg = 3'b111; end
            18'b100100100011101111: begin rgb_reg = 3'b111; end
            18'b100100100011110000: begin rgb_reg = 3'b111; end
            18'b100100100011110111: begin rgb_reg = 3'b111; end
            18'b100100100011111000: begin rgb_reg = 3'b111; end
            18'b100100100011111011: begin rgb_reg = 3'b111; end
            18'b100100100011111100: begin rgb_reg = 3'b111; end
            18'b100100100100000011: begin rgb_reg = 3'b111; end
            18'b100100100100000100: begin rgb_reg = 3'b111; end
            18'b100100100100000111: begin rgb_reg = 3'b111; end
            18'b100100100100001000: begin rgb_reg = 3'b111; end
            18'b100100100100001011: begin rgb_reg = 3'b111; end
            18'b100100100100001100: begin rgb_reg = 3'b111; end
            18'b100100100100001111: begin rgb_reg = 3'b111; end
            18'b100100100100010000: begin rgb_reg = 3'b111; end
            18'b100100100100010101: begin rgb_reg = 3'b111; end
            18'b100100100100010110: begin rgb_reg = 3'b111; end
            18'b100100100100010111: begin rgb_reg = 3'b111; end
            18'b100100100100011000: begin rgb_reg = 3'b111; end
            18'b100100100100011001: begin rgb_reg = 3'b111; end
            18'b100100100100011010: begin rgb_reg = 3'b111; end
            18'b100100100100011011: begin rgb_reg = 3'b111; end
            18'b100100100100011100: begin rgb_reg = 3'b111; end
            18'b100100100100011111: begin rgb_reg = 3'b111; end
            18'b100100100100100000: begin rgb_reg = 3'b111; end
            18'b100100100100100111: begin rgb_reg = 3'b111; end
            18'b100100100100101000: begin rgb_reg = 3'b111; end
            18'b100100100100101101: begin rgb_reg = 3'b111; end
            18'b100100100100101110: begin rgb_reg = 3'b111; end
            18'b100100100100101111: begin rgb_reg = 3'b111; end
            18'b100100100100110000: begin rgb_reg = 3'b111; end
            18'b100100100100110001: begin rgb_reg = 3'b111; end
            18'b100100100100110010: begin rgb_reg = 3'b111; end
            18'b100100100100110111: begin rgb_reg = 3'b111; end
            18'b100100100100111000: begin rgb_reg = 3'b111; end
            18'b100100100100111011: begin rgb_reg = 3'b111; end
            18'b100100100100111100: begin rgb_reg = 3'b111; end
            18'b100100100101000011: begin rgb_reg = 3'b111; end
            18'b100100100101000100: begin rgb_reg = 3'b111; end
            18'b100100100101000111: begin rgb_reg = 3'b111; end
            18'b100100100101001000: begin rgb_reg = 3'b111; end
            18'b100100100101001111: begin rgb_reg = 3'b111; end
            18'b100100100101010000: begin rgb_reg = 3'b111; end
            18'b100100100101010011: begin rgb_reg = 3'b111; end
            18'b100100100101010100: begin rgb_reg = 3'b111; end
            18'b100100100101011011: begin rgb_reg = 3'b111; end
            18'b100100100101011100: begin rgb_reg = 3'b111; end
            18'b100100100101100001: begin rgb_reg = 3'b111; end
            18'b100100100101100010: begin rgb_reg = 3'b111; end
            18'b100100100101100011: begin rgb_reg = 3'b111; end
            18'b100100100101100100: begin rgb_reg = 3'b111; end
            18'b100100100101100101: begin rgb_reg = 3'b111; end
            18'b100100100101100110: begin rgb_reg = 3'b111; end
            18'b100100100101100111: begin rgb_reg = 3'b111; end
            18'b100100100101101000: begin rgb_reg = 3'b111; end
            18'b100100100101101011: begin rgb_reg = 3'b111; end
            18'b100100100101101100: begin rgb_reg = 3'b111; end
            18'b100100100101110011: begin rgb_reg = 3'b111; end
            18'b100100100101110100: begin rgb_reg = 3'b111; end
            18'b100100100101111001: begin rgb_reg = 3'b111; end
            18'b100100100101111010: begin rgb_reg = 3'b111; end
            18'b100100100101111011: begin rgb_reg = 3'b111; end
            18'b100100100101111100: begin rgb_reg = 3'b111; end
            18'b100100100101111101: begin rgb_reg = 3'b111; end
            18'b100100100101111110: begin rgb_reg = 3'b111; end
            18'b100100100101111111: begin rgb_reg = 3'b111; end
            18'b100100100110000000: begin rgb_reg = 3'b111; end
            18'b100100100110000101: begin rgb_reg = 3'b111; end
            18'b100100100110000110: begin rgb_reg = 3'b111; end
            18'b100100101001111011: begin rgb_reg = 3'b111; end
            18'b100100101001111100: begin rgb_reg = 3'b111; end
            18'b100100101010000011: begin rgb_reg = 3'b111; end
            18'b100100101010000100: begin rgb_reg = 3'b111; end
            18'b100100101010001011: begin rgb_reg = 3'b111; end
            18'b100100101010001100: begin rgb_reg = 3'b111; end
            18'b100100101010001111: begin rgb_reg = 3'b111; end
            18'b100100101010010000: begin rgb_reg = 3'b111; end
            18'b100100101010010111: begin rgb_reg = 3'b111; end
            18'b100100101010011000: begin rgb_reg = 3'b111; end
            18'b100100101010011011: begin rgb_reg = 3'b111; end
            18'b100100101010011100: begin rgb_reg = 3'b111; end
            18'b100100101010011111: begin rgb_reg = 3'b111; end
            18'b100100101010100000: begin rgb_reg = 3'b111; end
            18'b100100101010100011: begin rgb_reg = 3'b111; end
            18'b100100101010100100: begin rgb_reg = 3'b111; end
            18'b100100101010100111: begin rgb_reg = 3'b111; end
            18'b100100101010101000: begin rgb_reg = 3'b111; end
            18'b100100101010101111: begin rgb_reg = 3'b111; end
            18'b100100101010110000: begin rgb_reg = 3'b111; end
            18'b100100101010110011: begin rgb_reg = 3'b111; end
            18'b100100101010110100: begin rgb_reg = 3'b111; end
            18'b100100101010111111: begin rgb_reg = 3'b111; end
            18'b100100101011000000: begin rgb_reg = 3'b111; end
            18'b100100101011000111: begin rgb_reg = 3'b111; end
            18'b100100101011001000: begin rgb_reg = 3'b111; end
            18'b100100101011010111: begin rgb_reg = 3'b111; end
            18'b100100101011011000: begin rgb_reg = 3'b111; end
            18'b100100101011011111: begin rgb_reg = 3'b111; end
            18'b100100101011100000: begin rgb_reg = 3'b111; end
            18'b100100101011100011: begin rgb_reg = 3'b111; end
            18'b100100101011100100: begin rgb_reg = 3'b111; end
            18'b100100101011101011: begin rgb_reg = 3'b111; end
            18'b100100101011101100: begin rgb_reg = 3'b111; end
            18'b100100101011101111: begin rgb_reg = 3'b111; end
            18'b100100101011110000: begin rgb_reg = 3'b111; end
            18'b100100101011110111: begin rgb_reg = 3'b111; end
            18'b100100101011111000: begin rgb_reg = 3'b111; end
            18'b100100101011111101: begin rgb_reg = 3'b111; end
            18'b100100101011111110: begin rgb_reg = 3'b111; end
            18'b100100101011111111: begin rgb_reg = 3'b111; end
            18'b100100101100000000: begin rgb_reg = 3'b111; end
            18'b100100101100000001: begin rgb_reg = 3'b111; end
            18'b100100101100000010: begin rgb_reg = 3'b111; end
            18'b100100101100000011: begin rgb_reg = 3'b111; end
            18'b100100101100000100: begin rgb_reg = 3'b111; end
            18'b100100101100000111: begin rgb_reg = 3'b111; end
            18'b100100101100001000: begin rgb_reg = 3'b111; end
            18'b100100101100001011: begin rgb_reg = 3'b111; end
            18'b100100101100001100: begin rgb_reg = 3'b111; end
            18'b100100101100001111: begin rgb_reg = 3'b111; end
            18'b100100101100010000: begin rgb_reg = 3'b111; end
            18'b100100101100010011: begin rgb_reg = 3'b111; end
            18'b100100101100010100: begin rgb_reg = 3'b111; end
            18'b100100101100011011: begin rgb_reg = 3'b111; end
            18'b100100101100011100: begin rgb_reg = 3'b111; end
            18'b100100101100011111: begin rgb_reg = 3'b111; end
            18'b100100101100100000: begin rgb_reg = 3'b111; end
            18'b100100101100100111: begin rgb_reg = 3'b111; end
            18'b100100101100101000: begin rgb_reg = 3'b111; end
            18'b100100101100110011: begin rgb_reg = 3'b111; end
            18'b100100101100110100: begin rgb_reg = 3'b111; end
            18'b100100101100110111: begin rgb_reg = 3'b111; end
            18'b100100101100111000: begin rgb_reg = 3'b111; end
            18'b100100101100111011: begin rgb_reg = 3'b111; end
            18'b100100101100111100: begin rgb_reg = 3'b111; end
            18'b100100101101000011: begin rgb_reg = 3'b111; end
            18'b100100101101000100: begin rgb_reg = 3'b111; end
            18'b100100101101001001: begin rgb_reg = 3'b111; end
            18'b100100101101001010: begin rgb_reg = 3'b111; end
            18'b100100101101001011: begin rgb_reg = 3'b111; end
            18'b100100101101001100: begin rgb_reg = 3'b111; end
            18'b100100101101001101: begin rgb_reg = 3'b111; end
            18'b100100101101001110: begin rgb_reg = 3'b111; end
            18'b100100101101001111: begin rgb_reg = 3'b111; end
            18'b100100101101010000: begin rgb_reg = 3'b111; end
            18'b100100101101010011: begin rgb_reg = 3'b111; end
            18'b100100101101010100: begin rgb_reg = 3'b111; end
            18'b100100101101011011: begin rgb_reg = 3'b111; end
            18'b100100101101011100: begin rgb_reg = 3'b111; end
            18'b100100101101011111: begin rgb_reg = 3'b111; end
            18'b100100101101100000: begin rgb_reg = 3'b111; end
            18'b100100101101100111: begin rgb_reg = 3'b111; end
            18'b100100101101101000: begin rgb_reg = 3'b111; end
            18'b100100101101101011: begin rgb_reg = 3'b111; end
            18'b100100101101101100: begin rgb_reg = 3'b111; end
            18'b100100101101110011: begin rgb_reg = 3'b111; end
            18'b100100101101110100: begin rgb_reg = 3'b111; end
            18'b100100101101110111: begin rgb_reg = 3'b111; end
            18'b100100101101111000: begin rgb_reg = 3'b111; end
            18'b100100101101111111: begin rgb_reg = 3'b111; end
            18'b100100101110000000: begin rgb_reg = 3'b111; end
            18'b100100101110000101: begin rgb_reg = 3'b111; end
            18'b100100101110000110: begin rgb_reg = 3'b111; end
            18'b100100110001111011: begin rgb_reg = 3'b111; end
            18'b100100110001111100: begin rgb_reg = 3'b111; end
            18'b100100110010000011: begin rgb_reg = 3'b111; end
            18'b100100110010000100: begin rgb_reg = 3'b111; end
            18'b100100110010001011: begin rgb_reg = 3'b111; end
            18'b100100110010001100: begin rgb_reg = 3'b111; end
            18'b100100110010001111: begin rgb_reg = 3'b111; end
            18'b100100110010010000: begin rgb_reg = 3'b111; end
            18'b100100110010010111: begin rgb_reg = 3'b111; end
            18'b100100110010011000: begin rgb_reg = 3'b111; end
            18'b100100110010011011: begin rgb_reg = 3'b111; end
            18'b100100110010011100: begin rgb_reg = 3'b111; end
            18'b100100110010011111: begin rgb_reg = 3'b111; end
            18'b100100110010100000: begin rgb_reg = 3'b111; end
            18'b100100110010100011: begin rgb_reg = 3'b111; end
            18'b100100110010100100: begin rgb_reg = 3'b111; end
            18'b100100110010100111: begin rgb_reg = 3'b111; end
            18'b100100110010101000: begin rgb_reg = 3'b111; end
            18'b100100110010101111: begin rgb_reg = 3'b111; end
            18'b100100110010110000: begin rgb_reg = 3'b111; end
            18'b100100110010110011: begin rgb_reg = 3'b111; end
            18'b100100110010110100: begin rgb_reg = 3'b111; end
            18'b100100110010111111: begin rgb_reg = 3'b111; end
            18'b100100110011000000: begin rgb_reg = 3'b111; end
            18'b100100110011000111: begin rgb_reg = 3'b111; end
            18'b100100110011001000: begin rgb_reg = 3'b111; end
            18'b100100110011010111: begin rgb_reg = 3'b111; end
            18'b100100110011011000: begin rgb_reg = 3'b111; end
            18'b100100110011011111: begin rgb_reg = 3'b111; end
            18'b100100110011100000: begin rgb_reg = 3'b111; end
            18'b100100110011100011: begin rgb_reg = 3'b111; end
            18'b100100110011100100: begin rgb_reg = 3'b111; end
            18'b100100110011101011: begin rgb_reg = 3'b111; end
            18'b100100110011101100: begin rgb_reg = 3'b111; end
            18'b100100110011101111: begin rgb_reg = 3'b111; end
            18'b100100110011110000: begin rgb_reg = 3'b111; end
            18'b100100110011110111: begin rgb_reg = 3'b111; end
            18'b100100110011111000: begin rgb_reg = 3'b111; end
            18'b100100110011111101: begin rgb_reg = 3'b111; end
            18'b100100110011111110: begin rgb_reg = 3'b111; end
            18'b100100110011111111: begin rgb_reg = 3'b111; end
            18'b100100110100000000: begin rgb_reg = 3'b111; end
            18'b100100110100000001: begin rgb_reg = 3'b111; end
            18'b100100110100000010: begin rgb_reg = 3'b111; end
            18'b100100110100000011: begin rgb_reg = 3'b111; end
            18'b100100110100000100: begin rgb_reg = 3'b111; end
            18'b100100110100000111: begin rgb_reg = 3'b111; end
            18'b100100110100001000: begin rgb_reg = 3'b111; end
            18'b100100110100001011: begin rgb_reg = 3'b111; end
            18'b100100110100001100: begin rgb_reg = 3'b111; end
            18'b100100110100001111: begin rgb_reg = 3'b111; end
            18'b100100110100010000: begin rgb_reg = 3'b111; end
            18'b100100110100010011: begin rgb_reg = 3'b111; end
            18'b100100110100010100: begin rgb_reg = 3'b111; end
            18'b100100110100011011: begin rgb_reg = 3'b111; end
            18'b100100110100011100: begin rgb_reg = 3'b111; end
            18'b100100110100011111: begin rgb_reg = 3'b111; end
            18'b100100110100100000: begin rgb_reg = 3'b111; end
            18'b100100110100100111: begin rgb_reg = 3'b111; end
            18'b100100110100101000: begin rgb_reg = 3'b111; end
            18'b100100110100110011: begin rgb_reg = 3'b111; end
            18'b100100110100110100: begin rgb_reg = 3'b111; end
            18'b100100110100110111: begin rgb_reg = 3'b111; end
            18'b100100110100111000: begin rgb_reg = 3'b111; end
            18'b100100110100111011: begin rgb_reg = 3'b111; end
            18'b100100110100111100: begin rgb_reg = 3'b111; end
            18'b100100110101000011: begin rgb_reg = 3'b111; end
            18'b100100110101000100: begin rgb_reg = 3'b111; end
            18'b100100110101001001: begin rgb_reg = 3'b111; end
            18'b100100110101001010: begin rgb_reg = 3'b111; end
            18'b100100110101001011: begin rgb_reg = 3'b111; end
            18'b100100110101001100: begin rgb_reg = 3'b111; end
            18'b100100110101001101: begin rgb_reg = 3'b111; end
            18'b100100110101001110: begin rgb_reg = 3'b111; end
            18'b100100110101001111: begin rgb_reg = 3'b111; end
            18'b100100110101010000: begin rgb_reg = 3'b111; end
            18'b100100110101010011: begin rgb_reg = 3'b111; end
            18'b100100110101010100: begin rgb_reg = 3'b111; end
            18'b100100110101011011: begin rgb_reg = 3'b111; end
            18'b100100110101011100: begin rgb_reg = 3'b111; end
            18'b100100110101011111: begin rgb_reg = 3'b111; end
            18'b100100110101100000: begin rgb_reg = 3'b111; end
            18'b100100110101100111: begin rgb_reg = 3'b111; end
            18'b100100110101101000: begin rgb_reg = 3'b111; end
            18'b100100110101101011: begin rgb_reg = 3'b111; end
            18'b100100110101101100: begin rgb_reg = 3'b111; end
            18'b100100110101110011: begin rgb_reg = 3'b111; end
            18'b100100110101110100: begin rgb_reg = 3'b111; end
            18'b100100110101110111: begin rgb_reg = 3'b111; end
            18'b100100110101111000: begin rgb_reg = 3'b111; end
            18'b100100110101111111: begin rgb_reg = 3'b111; end
            18'b100100110110000000: begin rgb_reg = 3'b111; end
            18'b100100110110000101: begin rgb_reg = 3'b111; end
            18'b100100110110000110: begin rgb_reg = 3'b111; end
            18'b100100111001111011: begin rgb_reg = 3'b111; end
            18'b100100111001111100: begin rgb_reg = 3'b111; end
            18'b100100111010000011: begin rgb_reg = 3'b111; end
            18'b100100111010000100: begin rgb_reg = 3'b111; end
            18'b100100111010001011: begin rgb_reg = 3'b111; end
            18'b100100111010001100: begin rgb_reg = 3'b111; end
            18'b100100111010010001: begin rgb_reg = 3'b111; end
            18'b100100111010010010: begin rgb_reg = 3'b111; end
            18'b100100111010010011: begin rgb_reg = 3'b111; end
            18'b100100111010010100: begin rgb_reg = 3'b111; end
            18'b100100111010010101: begin rgb_reg = 3'b111; end
            18'b100100111010010110: begin rgb_reg = 3'b111; end
            18'b100100111010010111: begin rgb_reg = 3'b111; end
            18'b100100111010011000: begin rgb_reg = 3'b111; end
            18'b100100111010011101: begin rgb_reg = 3'b111; end
            18'b100100111010011110: begin rgb_reg = 3'b111; end
            18'b100100111010011111: begin rgb_reg = 3'b111; end
            18'b100100111010100000: begin rgb_reg = 3'b111; end
            18'b100100111010100001: begin rgb_reg = 3'b111; end
            18'b100100111010100010: begin rgb_reg = 3'b111; end
            18'b100100111010100011: begin rgb_reg = 3'b111; end
            18'b100100111010100100: begin rgb_reg = 3'b111; end
            18'b100100111010101001: begin rgb_reg = 3'b111; end
            18'b100100111010101010: begin rgb_reg = 3'b111; end
            18'b100100111010101011: begin rgb_reg = 3'b111; end
            18'b100100111010101100: begin rgb_reg = 3'b111; end
            18'b100100111010101101: begin rgb_reg = 3'b111; end
            18'b100100111010101110: begin rgb_reg = 3'b111; end
            18'b100100111010110011: begin rgb_reg = 3'b111; end
            18'b100100111010110100: begin rgb_reg = 3'b111; end
            18'b100100111010111111: begin rgb_reg = 3'b111; end
            18'b100100111011000000: begin rgb_reg = 3'b111; end
            18'b100100111011000111: begin rgb_reg = 3'b111; end
            18'b100100111011001000: begin rgb_reg = 3'b111; end
            18'b100100111011010111: begin rgb_reg = 3'b111; end
            18'b100100111011011000: begin rgb_reg = 3'b111; end
            18'b100100111011011111: begin rgb_reg = 3'b111; end
            18'b100100111011100000: begin rgb_reg = 3'b111; end
            18'b100100111011100101: begin rgb_reg = 3'b111; end
            18'b100100111011100110: begin rgb_reg = 3'b111; end
            18'b100100111011100111: begin rgb_reg = 3'b111; end
            18'b100100111011101000: begin rgb_reg = 3'b111; end
            18'b100100111011101001: begin rgb_reg = 3'b111; end
            18'b100100111011101010: begin rgb_reg = 3'b111; end
            18'b100100111011101011: begin rgb_reg = 3'b111; end
            18'b100100111011101100: begin rgb_reg = 3'b111; end
            18'b100100111011101111: begin rgb_reg = 3'b111; end
            18'b100100111011110000: begin rgb_reg = 3'b111; end
            18'b100100111011110111: begin rgb_reg = 3'b111; end
            18'b100100111011111000: begin rgb_reg = 3'b111; end
            18'b100100111100000011: begin rgb_reg = 3'b111; end
            18'b100100111100000100: begin rgb_reg = 3'b111; end
            18'b100100111100001001: begin rgb_reg = 3'b111; end
            18'b100100111100001010: begin rgb_reg = 3'b111; end
            18'b100100111100001011: begin rgb_reg = 3'b111; end
            18'b100100111100001100: begin rgb_reg = 3'b111; end
            18'b100100111100001101: begin rgb_reg = 3'b111; end
            18'b100100111100001110: begin rgb_reg = 3'b111; end
            18'b100100111100001111: begin rgb_reg = 3'b111; end
            18'b100100111100010000: begin rgb_reg = 3'b111; end
            18'b100100111100010101: begin rgb_reg = 3'b111; end
            18'b100100111100010110: begin rgb_reg = 3'b111; end
            18'b100100111100010111: begin rgb_reg = 3'b111; end
            18'b100100111100011000: begin rgb_reg = 3'b111; end
            18'b100100111100011001: begin rgb_reg = 3'b111; end
            18'b100100111100011010: begin rgb_reg = 3'b111; end
            18'b100100111100011011: begin rgb_reg = 3'b111; end
            18'b100100111100011100: begin rgb_reg = 3'b111; end
            18'b100100111100011111: begin rgb_reg = 3'b111; end
            18'b100100111100100000: begin rgb_reg = 3'b111; end
            18'b100100111100100111: begin rgb_reg = 3'b111; end
            18'b100100111100101000: begin rgb_reg = 3'b111; end
            18'b100100111100101011: begin rgb_reg = 3'b111; end
            18'b100100111100101100: begin rgb_reg = 3'b111; end
            18'b100100111100101101: begin rgb_reg = 3'b111; end
            18'b100100111100101110: begin rgb_reg = 3'b111; end
            18'b100100111100101111: begin rgb_reg = 3'b111; end
            18'b100100111100110000: begin rgb_reg = 3'b111; end
            18'b100100111100110001: begin rgb_reg = 3'b111; end
            18'b100100111100110010: begin rgb_reg = 3'b111; end
            18'b100100111100110111: begin rgb_reg = 3'b111; end
            18'b100100111100111000: begin rgb_reg = 3'b111; end
            18'b100100111100111011: begin rgb_reg = 3'b111; end
            18'b100100111100111100: begin rgb_reg = 3'b111; end
            18'b100100111101000011: begin rgb_reg = 3'b111; end
            18'b100100111101000100: begin rgb_reg = 3'b111; end
            18'b100100111101001111: begin rgb_reg = 3'b111; end
            18'b100100111101010000: begin rgb_reg = 3'b111; end
            18'b100100111101010011: begin rgb_reg = 3'b111; end
            18'b100100111101010100: begin rgb_reg = 3'b111; end
            18'b100100111101011011: begin rgb_reg = 3'b111; end
            18'b100100111101011100: begin rgb_reg = 3'b111; end
            18'b100100111101100001: begin rgb_reg = 3'b111; end
            18'b100100111101100010: begin rgb_reg = 3'b111; end
            18'b100100111101100011: begin rgb_reg = 3'b111; end
            18'b100100111101100100: begin rgb_reg = 3'b111; end
            18'b100100111101100101: begin rgb_reg = 3'b111; end
            18'b100100111101100110: begin rgb_reg = 3'b111; end
            18'b100100111101100111: begin rgb_reg = 3'b111; end
            18'b100100111101101000: begin rgb_reg = 3'b111; end
            18'b100100111101101011: begin rgb_reg = 3'b111; end
            18'b100100111101101100: begin rgb_reg = 3'b111; end
            18'b100100111101110011: begin rgb_reg = 3'b111; end
            18'b100100111101110100: begin rgb_reg = 3'b111; end
            18'b100100111101111001: begin rgb_reg = 3'b111; end
            18'b100100111101111010: begin rgb_reg = 3'b111; end
            18'b100100111101111011: begin rgb_reg = 3'b111; end
            18'b100100111101111100: begin rgb_reg = 3'b111; end
            18'b100100111101111101: begin rgb_reg = 3'b111; end
            18'b100100111101111110: begin rgb_reg = 3'b111; end
            18'b100100111101111111: begin rgb_reg = 3'b111; end
            18'b100100111110000000: begin rgb_reg = 3'b111; end
            18'b100100111110000111: begin rgb_reg = 3'b111; end
            18'b100100111110001000: begin rgb_reg = 3'b111; end
            18'b100101000001111011: begin rgb_reg = 3'b111; end
            18'b100101000001111100: begin rgb_reg = 3'b111; end
            18'b100101000010000011: begin rgb_reg = 3'b111; end
            18'b100101000010000100: begin rgb_reg = 3'b111; end
            18'b100101000010001011: begin rgb_reg = 3'b111; end
            18'b100101000010001100: begin rgb_reg = 3'b111; end
            18'b100101000010010001: begin rgb_reg = 3'b111; end
            18'b100101000010010010: begin rgb_reg = 3'b111; end
            18'b100101000010010011: begin rgb_reg = 3'b111; end
            18'b100101000010010100: begin rgb_reg = 3'b111; end
            18'b100101000010010101: begin rgb_reg = 3'b111; end
            18'b100101000010010110: begin rgb_reg = 3'b111; end
            18'b100101000010010111: begin rgb_reg = 3'b111; end
            18'b100101000010011000: begin rgb_reg = 3'b111; end
            18'b100101000010011101: begin rgb_reg = 3'b111; end
            18'b100101000010011110: begin rgb_reg = 3'b111; end
            18'b100101000010011111: begin rgb_reg = 3'b111; end
            18'b100101000010100000: begin rgb_reg = 3'b111; end
            18'b100101000010100001: begin rgb_reg = 3'b111; end
            18'b100101000010100010: begin rgb_reg = 3'b111; end
            18'b100101000010100011: begin rgb_reg = 3'b111; end
            18'b100101000010100100: begin rgb_reg = 3'b111; end
            18'b100101000010101001: begin rgb_reg = 3'b111; end
            18'b100101000010101010: begin rgb_reg = 3'b111; end
            18'b100101000010101011: begin rgb_reg = 3'b111; end
            18'b100101000010101100: begin rgb_reg = 3'b111; end
            18'b100101000010101101: begin rgb_reg = 3'b111; end
            18'b100101000010101110: begin rgb_reg = 3'b111; end
            18'b100101000010110011: begin rgb_reg = 3'b111; end
            18'b100101000010110100: begin rgb_reg = 3'b111; end
            18'b100101000010111111: begin rgb_reg = 3'b111; end
            18'b100101000011000000: begin rgb_reg = 3'b111; end
            18'b100101000011000111: begin rgb_reg = 3'b111; end
            18'b100101000011001000: begin rgb_reg = 3'b111; end
            18'b100101000011010111: begin rgb_reg = 3'b111; end
            18'b100101000011011000: begin rgb_reg = 3'b111; end
            18'b100101000011011111: begin rgb_reg = 3'b111; end
            18'b100101000011100000: begin rgb_reg = 3'b111; end
            18'b100101000011100101: begin rgb_reg = 3'b111; end
            18'b100101000011100110: begin rgb_reg = 3'b111; end
            18'b100101000011100111: begin rgb_reg = 3'b111; end
            18'b100101000011101000: begin rgb_reg = 3'b111; end
            18'b100101000011101001: begin rgb_reg = 3'b111; end
            18'b100101000011101010: begin rgb_reg = 3'b111; end
            18'b100101000011101011: begin rgb_reg = 3'b111; end
            18'b100101000011101100: begin rgb_reg = 3'b111; end
            18'b100101000011101111: begin rgb_reg = 3'b111; end
            18'b100101000011110000: begin rgb_reg = 3'b111; end
            18'b100101000011110111: begin rgb_reg = 3'b111; end
            18'b100101000011111000: begin rgb_reg = 3'b111; end
            18'b100101000100000011: begin rgb_reg = 3'b111; end
            18'b100101000100000100: begin rgb_reg = 3'b111; end
            18'b100101000100001001: begin rgb_reg = 3'b111; end
            18'b100101000100001010: begin rgb_reg = 3'b111; end
            18'b100101000100001011: begin rgb_reg = 3'b111; end
            18'b100101000100001100: begin rgb_reg = 3'b111; end
            18'b100101000100001101: begin rgb_reg = 3'b111; end
            18'b100101000100001110: begin rgb_reg = 3'b111; end
            18'b100101000100001111: begin rgb_reg = 3'b111; end
            18'b100101000100010000: begin rgb_reg = 3'b111; end
            18'b100101000100010101: begin rgb_reg = 3'b111; end
            18'b100101000100010110: begin rgb_reg = 3'b111; end
            18'b100101000100010111: begin rgb_reg = 3'b111; end
            18'b100101000100011000: begin rgb_reg = 3'b111; end
            18'b100101000100011001: begin rgb_reg = 3'b111; end
            18'b100101000100011010: begin rgb_reg = 3'b111; end
            18'b100101000100011011: begin rgb_reg = 3'b111; end
            18'b100101000100011100: begin rgb_reg = 3'b111; end
            18'b100101000100011111: begin rgb_reg = 3'b111; end
            18'b100101000100100000: begin rgb_reg = 3'b111; end
            18'b100101000100100111: begin rgb_reg = 3'b111; end
            18'b100101000100101000: begin rgb_reg = 3'b111; end
            18'b100101000100101011: begin rgb_reg = 3'b111; end
            18'b100101000100101100: begin rgb_reg = 3'b111; end
            18'b100101000100101101: begin rgb_reg = 3'b111; end
            18'b100101000100101110: begin rgb_reg = 3'b111; end
            18'b100101000100101111: begin rgb_reg = 3'b111; end
            18'b100101000100110000: begin rgb_reg = 3'b111; end
            18'b100101000100110001: begin rgb_reg = 3'b111; end
            18'b100101000100110010: begin rgb_reg = 3'b111; end
            18'b100101000100110111: begin rgb_reg = 3'b111; end
            18'b100101000100111000: begin rgb_reg = 3'b111; end
            18'b100101000100111011: begin rgb_reg = 3'b111; end
            18'b100101000100111100: begin rgb_reg = 3'b111; end
            18'b100101000101000011: begin rgb_reg = 3'b111; end
            18'b100101000101000100: begin rgb_reg = 3'b111; end
            18'b100101000101001111: begin rgb_reg = 3'b111; end
            18'b100101000101010000: begin rgb_reg = 3'b111; end
            18'b100101000101010011: begin rgb_reg = 3'b111; end
            18'b100101000101010100: begin rgb_reg = 3'b111; end
            18'b100101000101011011: begin rgb_reg = 3'b111; end
            18'b100101000101011100: begin rgb_reg = 3'b111; end
            18'b100101000101100001: begin rgb_reg = 3'b111; end
            18'b100101000101100010: begin rgb_reg = 3'b111; end
            18'b100101000101100011: begin rgb_reg = 3'b111; end
            18'b100101000101100100: begin rgb_reg = 3'b111; end
            18'b100101000101100101: begin rgb_reg = 3'b111; end
            18'b100101000101100110: begin rgb_reg = 3'b111; end
            18'b100101000101100111: begin rgb_reg = 3'b111; end
            18'b100101000101101000: begin rgb_reg = 3'b111; end
            18'b100101000101101011: begin rgb_reg = 3'b111; end
            18'b100101000101101100: begin rgb_reg = 3'b111; end
            18'b100101000101110011: begin rgb_reg = 3'b111; end
            18'b100101000101110100: begin rgb_reg = 3'b111; end
            18'b100101000101111001: begin rgb_reg = 3'b111; end
            18'b100101000101111010: begin rgb_reg = 3'b111; end
            18'b100101000101111011: begin rgb_reg = 3'b111; end
            18'b100101000101111100: begin rgb_reg = 3'b111; end
            18'b100101000101111101: begin rgb_reg = 3'b111; end
            18'b100101000101111110: begin rgb_reg = 3'b111; end
            18'b100101000101111111: begin rgb_reg = 3'b111; end
            18'b100101000110000000: begin rgb_reg = 3'b111; end
            18'b100101000110000111: begin rgb_reg = 3'b111; end
            18'b100101000110001000: begin rgb_reg = 3'b111; end
            18'b100101001011111011: begin rgb_reg = 3'b111; end
            18'b100101001011111100: begin rgb_reg = 3'b111; end
            18'b100101001011111101: begin rgb_reg = 3'b111; end
            18'b100101001011111110: begin rgb_reg = 3'b111; end
            18'b100101001011111111: begin rgb_reg = 3'b111; end
            18'b100101001100000000: begin rgb_reg = 3'b111; end
            18'b100101001100000001: begin rgb_reg = 3'b111; end
            18'b100101001100000010: begin rgb_reg = 3'b111; end
            18'b100101001101000111: begin rgb_reg = 3'b111; end
            18'b100101001101001000: begin rgb_reg = 3'b111; end
            18'b100101001101001001: begin rgb_reg = 3'b111; end
            18'b100101001101001010: begin rgb_reg = 3'b111; end
            18'b100101001101001011: begin rgb_reg = 3'b111; end
            18'b100101001101001100: begin rgb_reg = 3'b111; end
            18'b100101001101001101: begin rgb_reg = 3'b111; end
            18'b100101001101001110: begin rgb_reg = 3'b111; end
            18'b100101010011111011: begin rgb_reg = 3'b111; end
            18'b100101010011111100: begin rgb_reg = 3'b111; end
            18'b100101010011111101: begin rgb_reg = 3'b111; end
            18'b100101010011111110: begin rgb_reg = 3'b111; end
            18'b100101010011111111: begin rgb_reg = 3'b111; end
            18'b100101010100000000: begin rgb_reg = 3'b111; end
            18'b100101010100000001: begin rgb_reg = 3'b111; end
            18'b100101010100000010: begin rgb_reg = 3'b111; end
            18'b100101010101000111: begin rgb_reg = 3'b111; end
            18'b100101010101001000: begin rgb_reg = 3'b111; end
            18'b100101010101001001: begin rgb_reg = 3'b111; end
            18'b100101010101001010: begin rgb_reg = 3'b111; end
            18'b100101010101001011: begin rgb_reg = 3'b111; end
            18'b100101010101001100: begin rgb_reg = 3'b111; end
            18'b100101010101001101: begin rgb_reg = 3'b111; end
            18'b100101010101001110: begin rgb_reg = 3'b111; end
            18'b100111111011000010: begin rgb_reg = 3'b111; end
            18'b100111111011000011: begin rgb_reg = 3'b111; end
            18'b100111111011000100: begin rgb_reg = 3'b111; end
            18'b100111111011000101: begin rgb_reg = 3'b111; end
            18'b100111111011000110: begin rgb_reg = 3'b111; end
            18'b100111111011001101: begin rgb_reg = 3'b111; end
            18'b100111111011001110: begin rgb_reg = 3'b111; end
            18'b100111111011001111: begin rgb_reg = 3'b111; end
            18'b100111111011010000: begin rgb_reg = 3'b111; end
            18'b100111111011010001: begin rgb_reg = 3'b111; end
            18'b100111111011010010: begin rgb_reg = 3'b111; end
            18'b100111111011010011: begin rgb_reg = 3'b111; end
            18'b100111111011011011: begin rgb_reg = 3'b111; end
            18'b100111111011011100: begin rgb_reg = 3'b111; end
            18'b100111111011011101: begin rgb_reg = 3'b111; end
            18'b100111111011011110: begin rgb_reg = 3'b111; end
            18'b100111111011011111: begin rgb_reg = 3'b111; end
            18'b100111111011100000: begin rgb_reg = 3'b111; end
            18'b100111111011100001: begin rgb_reg = 3'b111; end
            18'b100111111011101011: begin rgb_reg = 3'b111; end
            18'b100111111011101100: begin rgb_reg = 3'b111; end
            18'b100111111011110110: begin rgb_reg = 3'b111; end
            18'b100111111011110111: begin rgb_reg = 3'b111; end
            18'b100111111011111000: begin rgb_reg = 3'b111; end
            18'b100111111011111001: begin rgb_reg = 3'b111; end
            18'b100111111011111010: begin rgb_reg = 3'b111; end
            18'b100111111011111011: begin rgb_reg = 3'b111; end
            18'b100111111011111100: begin rgb_reg = 3'b111; end
            18'b100111111100000110: begin rgb_reg = 3'b111; end
            18'b100111111100000111: begin rgb_reg = 3'b111; end
            18'b100111111100010101: begin rgb_reg = 3'b111; end
            18'b100111111100010110: begin rgb_reg = 3'b111; end
            18'b100111111100010111: begin rgb_reg = 3'b111; end
            18'b100111111100011000: begin rgb_reg = 3'b111; end
            18'b100111111100011001: begin rgb_reg = 3'b111; end
            18'b100111111100100001: begin rgb_reg = 3'b111; end
            18'b100111111100100010: begin rgb_reg = 3'b111; end
            18'b100111111100100011: begin rgb_reg = 3'b111; end
            18'b100111111100100100: begin rgb_reg = 3'b111; end
            18'b100111111100101100: begin rgb_reg = 3'b111; end
            18'b100111111100101101: begin rgb_reg = 3'b111; end
            18'b100111111100101110: begin rgb_reg = 3'b111; end
            18'b100111111100101111: begin rgb_reg = 3'b111; end
            18'b100111111100110000: begin rgb_reg = 3'b111; end
            18'b100111111100110001: begin rgb_reg = 3'b111; end
            18'b100111111100110010: begin rgb_reg = 3'b111; end
            18'b100111111100111100: begin rgb_reg = 3'b111; end
            18'b100111111100111101: begin rgb_reg = 3'b111; end
            18'b101000000011000010: begin rgb_reg = 3'b111; end
            18'b101000000011000011: begin rgb_reg = 3'b111; end
            18'b101000000011000100: begin rgb_reg = 3'b111; end
            18'b101000000011000101: begin rgb_reg = 3'b111; end
            18'b101000000011000110: begin rgb_reg = 3'b111; end
            18'b101000000011001101: begin rgb_reg = 3'b111; end
            18'b101000000011001110: begin rgb_reg = 3'b111; end
            18'b101000000011001111: begin rgb_reg = 3'b111; end
            18'b101000000011010000: begin rgb_reg = 3'b111; end
            18'b101000000011010001: begin rgb_reg = 3'b111; end
            18'b101000000011010010: begin rgb_reg = 3'b111; end
            18'b101000000011010011: begin rgb_reg = 3'b111; end
            18'b101000000011011011: begin rgb_reg = 3'b111; end
            18'b101000000011011100: begin rgb_reg = 3'b111; end
            18'b101000000011011101: begin rgb_reg = 3'b111; end
            18'b101000000011011110: begin rgb_reg = 3'b111; end
            18'b101000000011011111: begin rgb_reg = 3'b111; end
            18'b101000000011100000: begin rgb_reg = 3'b111; end
            18'b101000000011100001: begin rgb_reg = 3'b111; end
            18'b101000000011101011: begin rgb_reg = 3'b111; end
            18'b101000000011101100: begin rgb_reg = 3'b111; end
            18'b101000000011110110: begin rgb_reg = 3'b111; end
            18'b101000000011110111: begin rgb_reg = 3'b111; end
            18'b101000000011111000: begin rgb_reg = 3'b111; end
            18'b101000000011111001: begin rgb_reg = 3'b111; end
            18'b101000000011111010: begin rgb_reg = 3'b111; end
            18'b101000000011111011: begin rgb_reg = 3'b111; end
            18'b101000000011111100: begin rgb_reg = 3'b111; end
            18'b101000000100000110: begin rgb_reg = 3'b111; end
            18'b101000000100000111: begin rgb_reg = 3'b111; end
            18'b101000000100010101: begin rgb_reg = 3'b111; end
            18'b101000000100010110: begin rgb_reg = 3'b111; end
            18'b101000000100010111: begin rgb_reg = 3'b111; end
            18'b101000000100011000: begin rgb_reg = 3'b111; end
            18'b101000000100011001: begin rgb_reg = 3'b111; end
            18'b101000000100100001: begin rgb_reg = 3'b111; end
            18'b101000000100100010: begin rgb_reg = 3'b111; end
            18'b101000000100100011: begin rgb_reg = 3'b111; end
            18'b101000000100100100: begin rgb_reg = 3'b111; end
            18'b101000000100101100: begin rgb_reg = 3'b111; end
            18'b101000000100101101: begin rgb_reg = 3'b111; end
            18'b101000000100101110: begin rgb_reg = 3'b111; end
            18'b101000000100101111: begin rgb_reg = 3'b111; end
            18'b101000000100110000: begin rgb_reg = 3'b111; end
            18'b101000000100110001: begin rgb_reg = 3'b111; end
            18'b101000000100110010: begin rgb_reg = 3'b111; end
            18'b101000000100111100: begin rgb_reg = 3'b111; end
            18'b101000000100111101: begin rgb_reg = 3'b111; end
            18'b101000001011000000: begin rgb_reg = 3'b111; end
            18'b101000001011000001: begin rgb_reg = 3'b111; end
            18'b101000001011001011: begin rgb_reg = 3'b111; end
            18'b101000001011001100: begin rgb_reg = 3'b111; end
            18'b101000001011001101: begin rgb_reg = 3'b111; end
            18'b101000001011010100: begin rgb_reg = 3'b111; end
            18'b101000001011010101: begin rgb_reg = 3'b111; end
            18'b101000001011011001: begin rgb_reg = 3'b111; end
            18'b101000001011011010: begin rgb_reg = 3'b111; end
            18'b101000001011100010: begin rgb_reg = 3'b111; end
            18'b101000001011100011: begin rgb_reg = 3'b111; end
            18'b101000001011101001: begin rgb_reg = 3'b111; end
            18'b101000001011101010: begin rgb_reg = 3'b111; end
            18'b101000001011101011: begin rgb_reg = 3'b111; end
            18'b101000001011101100: begin rgb_reg = 3'b111; end
            18'b101000001011110100: begin rgb_reg = 3'b111; end
            18'b101000001011110101: begin rgb_reg = 3'b111; end
            18'b101000001011111101: begin rgb_reg = 3'b111; end
            18'b101000001011111110: begin rgb_reg = 3'b111; end
            18'b101000001100000100: begin rgb_reg = 3'b111; end
            18'b101000001100000101: begin rgb_reg = 3'b111; end
            18'b101000001100000110: begin rgb_reg = 3'b111; end
            18'b101000001100000111: begin rgb_reg = 3'b111; end
            18'b101000001100010011: begin rgb_reg = 3'b111; end
            18'b101000001100010100: begin rgb_reg = 3'b111; end
            18'b101000001100010101: begin rgb_reg = 3'b111; end
            18'b101000001100010111: begin rgb_reg = 3'b111; end
            18'b101000001100011000: begin rgb_reg = 3'b111; end
            18'b101000001100011001: begin rgb_reg = 3'b111; end
            18'b101000001100011111: begin rgb_reg = 3'b111; end
            18'b101000001100100000: begin rgb_reg = 3'b111; end
            18'b101000001100101010: begin rgb_reg = 3'b111; end
            18'b101000001100101011: begin rgb_reg = 3'b111; end
            18'b101000001100110011: begin rgb_reg = 3'b111; end
            18'b101000001100110100: begin rgb_reg = 3'b111; end
            18'b101000001100111010: begin rgb_reg = 3'b111; end
            18'b101000001100111011: begin rgb_reg = 3'b111; end
            18'b101000001100111100: begin rgb_reg = 3'b111; end
            18'b101000001100111101: begin rgb_reg = 3'b111; end
            18'b101000010011000000: begin rgb_reg = 3'b111; end
            18'b101000010011000001: begin rgb_reg = 3'b111; end
            18'b101000010011001011: begin rgb_reg = 3'b111; end
            18'b101000010011001100: begin rgb_reg = 3'b111; end
            18'b101000010011001101: begin rgb_reg = 3'b111; end
            18'b101000010011010100: begin rgb_reg = 3'b111; end
            18'b101000010011010101: begin rgb_reg = 3'b111; end
            18'b101000010011010110: begin rgb_reg = 3'b111; end
            18'b101000010011011001: begin rgb_reg = 3'b111; end
            18'b101000010011011010: begin rgb_reg = 3'b111; end
            18'b101000010011100010: begin rgb_reg = 3'b111; end
            18'b101000010011100011: begin rgb_reg = 3'b111; end
            18'b101000010011101000: begin rgb_reg = 3'b111; end
            18'b101000010011101001: begin rgb_reg = 3'b111; end
            18'b101000010011101010: begin rgb_reg = 3'b111; end
            18'b101000010011101011: begin rgb_reg = 3'b111; end
            18'b101000010011101100: begin rgb_reg = 3'b111; end
            18'b101000010011110100: begin rgb_reg = 3'b111; end
            18'b101000010011110101: begin rgb_reg = 3'b111; end
            18'b101000010011111101: begin rgb_reg = 3'b111; end
            18'b101000010011111110: begin rgb_reg = 3'b111; end
            18'b101000010100000011: begin rgb_reg = 3'b111; end
            18'b101000010100000100: begin rgb_reg = 3'b111; end
            18'b101000010100000101: begin rgb_reg = 3'b111; end
            18'b101000010100000110: begin rgb_reg = 3'b111; end
            18'b101000010100000111: begin rgb_reg = 3'b111; end
            18'b101000010100010011: begin rgb_reg = 3'b111; end
            18'b101000010100010100: begin rgb_reg = 3'b111; end
            18'b101000010100010101: begin rgb_reg = 3'b111; end
            18'b101000010100011000: begin rgb_reg = 3'b111; end
            18'b101000010100011001: begin rgb_reg = 3'b111; end
            18'b101000010100011110: begin rgb_reg = 3'b111; end
            18'b101000010100011111: begin rgb_reg = 3'b111; end
            18'b101000010100100000: begin rgb_reg = 3'b111; end
            18'b101000010100101010: begin rgb_reg = 3'b111; end
            18'b101000010100101011: begin rgb_reg = 3'b111; end
            18'b101000010100110011: begin rgb_reg = 3'b111; end
            18'b101000010100110100: begin rgb_reg = 3'b111; end
            18'b101000010100111001: begin rgb_reg = 3'b111; end
            18'b101000010100111010: begin rgb_reg = 3'b111; end
            18'b101000010100111011: begin rgb_reg = 3'b111; end
            18'b101000010100111100: begin rgb_reg = 3'b111; end
            18'b101000010100111101: begin rgb_reg = 3'b111; end
            18'b101000011010111110: begin rgb_reg = 3'b111; end
            18'b101000011010111111: begin rgb_reg = 3'b111; end
            18'b101000011011000000: begin rgb_reg = 3'b111; end
            18'b101000011011000001: begin rgb_reg = 3'b111; end
            18'b101000011011001011: begin rgb_reg = 3'b111; end
            18'b101000011011001100: begin rgb_reg = 3'b111; end
            18'b101000011011001101: begin rgb_reg = 3'b111; end
            18'b101000011011010010: begin rgb_reg = 3'b111; end
            18'b101000011011010011: begin rgb_reg = 3'b111; end
            18'b101000011011010100: begin rgb_reg = 3'b111; end
            18'b101000011011010101: begin rgb_reg = 3'b111; end
            18'b101000011011010110: begin rgb_reg = 3'b111; end
            18'b101000011011011001: begin rgb_reg = 3'b111; end
            18'b101000011011011010: begin rgb_reg = 3'b111; end
            18'b101000011011100010: begin rgb_reg = 3'b111; end
            18'b101000011011100011: begin rgb_reg = 3'b111; end
            18'b101000011011101001: begin rgb_reg = 3'b111; end
            18'b101000011011101010: begin rgb_reg = 3'b111; end
            18'b101000011011101011: begin rgb_reg = 3'b111; end
            18'b101000011011101100: begin rgb_reg = 3'b111; end
            18'b101000011011110100: begin rgb_reg = 3'b111; end
            18'b101000011011110101: begin rgb_reg = 3'b111; end
            18'b101000011011111011: begin rgb_reg = 3'b111; end
            18'b101000011011111100: begin rgb_reg = 3'b111; end
            18'b101000011011111101: begin rgb_reg = 3'b111; end
            18'b101000011011111110: begin rgb_reg = 3'b111; end
            18'b101000011100000100: begin rgb_reg = 3'b111; end
            18'b101000011100000101: begin rgb_reg = 3'b111; end
            18'b101000011100000110: begin rgb_reg = 3'b111; end
            18'b101000011100000111: begin rgb_reg = 3'b111; end
            18'b101000011100010001: begin rgb_reg = 3'b111; end
            18'b101000011100010010: begin rgb_reg = 3'b111; end
            18'b101000011100010011: begin rgb_reg = 3'b111; end
            18'b101000011100010100: begin rgb_reg = 3'b111; end
            18'b101000011100011000: begin rgb_reg = 3'b111; end
            18'b101000011100011001: begin rgb_reg = 3'b111; end
            18'b101000011100011101: begin rgb_reg = 3'b111; end
            18'b101000011100011110: begin rgb_reg = 3'b111; end
            18'b101000011100011111: begin rgb_reg = 3'b111; end
            18'b101000011100101010: begin rgb_reg = 3'b111; end
            18'b101000011100101011: begin rgb_reg = 3'b111; end
            18'b101000011100110011: begin rgb_reg = 3'b111; end
            18'b101000011100110100: begin rgb_reg = 3'b111; end
            18'b101000011100111010: begin rgb_reg = 3'b111; end
            18'b101000011100111011: begin rgb_reg = 3'b111; end
            18'b101000011100111100: begin rgb_reg = 3'b111; end
            18'b101000011100111101: begin rgb_reg = 3'b111; end
            18'b101000100010111110: begin rgb_reg = 3'b111; end
            18'b101000100010111111: begin rgb_reg = 3'b111; end
            18'b101000100011001011: begin rgb_reg = 3'b111; end
            18'b101000100011001100: begin rgb_reg = 3'b111; end
            18'b101000100011001101: begin rgb_reg = 3'b111; end
            18'b101000100011010010: begin rgb_reg = 3'b111; end
            18'b101000100011010011: begin rgb_reg = 3'b111; end
            18'b101000100011010100: begin rgb_reg = 3'b111; end
            18'b101000100011010101: begin rgb_reg = 3'b111; end
            18'b101000100011010110: begin rgb_reg = 3'b111; end
            18'b101000100011100010: begin rgb_reg = 3'b111; end
            18'b101000100011100011: begin rgb_reg = 3'b111; end
            18'b101000100011101011: begin rgb_reg = 3'b111; end
            18'b101000100011101100: begin rgb_reg = 3'b111; end
            18'b101000100011110100: begin rgb_reg = 3'b111; end
            18'b101000100011110101: begin rgb_reg = 3'b111; end
            18'b101000100011111010: begin rgb_reg = 3'b111; end
            18'b101000100011111011: begin rgb_reg = 3'b111; end
            18'b101000100011111100: begin rgb_reg = 3'b111; end
            18'b101000100011111101: begin rgb_reg = 3'b111; end
            18'b101000100011111110: begin rgb_reg = 3'b111; end
            18'b101000100100000110: begin rgb_reg = 3'b111; end
            18'b101000100100000111: begin rgb_reg = 3'b111; end
            18'b101000100100010001: begin rgb_reg = 3'b111; end
            18'b101000100100010010: begin rgb_reg = 3'b111; end
            18'b101000100100011000: begin rgb_reg = 3'b111; end
            18'b101000100100011001: begin rgb_reg = 3'b111; end
            18'b101000100100011100: begin rgb_reg = 3'b111; end
            18'b101000100100011101: begin rgb_reg = 3'b111; end
            18'b101000100100011110: begin rgb_reg = 3'b111; end
            18'b101000100100110011: begin rgb_reg = 3'b111; end
            18'b101000100100110100: begin rgb_reg = 3'b111; end
            18'b101000100100111100: begin rgb_reg = 3'b111; end
            18'b101000100100111101: begin rgb_reg = 3'b111; end
            18'b101000101010111110: begin rgb_reg = 3'b111; end
            18'b101000101010111111: begin rgb_reg = 3'b111; end
            18'b101000101011001011: begin rgb_reg = 3'b111; end
            18'b101000101011001100: begin rgb_reg = 3'b111; end
            18'b101000101011001101: begin rgb_reg = 3'b111; end
            18'b101000101011010010: begin rgb_reg = 3'b111; end
            18'b101000101011010011: begin rgb_reg = 3'b111; end
            18'b101000101011010100: begin rgb_reg = 3'b111; end
            18'b101000101011010101: begin rgb_reg = 3'b111; end
            18'b101000101011010110: begin rgb_reg = 3'b111; end
            18'b101000101011100010: begin rgb_reg = 3'b111; end
            18'b101000101011100011: begin rgb_reg = 3'b111; end
            18'b101000101011101011: begin rgb_reg = 3'b111; end
            18'b101000101011101100: begin rgb_reg = 3'b111; end
            18'b101000101011110100: begin rgb_reg = 3'b111; end
            18'b101000101011110101: begin rgb_reg = 3'b111; end
            18'b101000101011111010: begin rgb_reg = 3'b111; end
            18'b101000101011111011: begin rgb_reg = 3'b111; end
            18'b101000101011111100: begin rgb_reg = 3'b111; end
            18'b101000101011111101: begin rgb_reg = 3'b111; end
            18'b101000101011111110: begin rgb_reg = 3'b111; end
            18'b101000101100000110: begin rgb_reg = 3'b111; end
            18'b101000101100000111: begin rgb_reg = 3'b111; end
            18'b101000101100010001: begin rgb_reg = 3'b111; end
            18'b101000101100010010: begin rgb_reg = 3'b111; end
            18'b101000101100011000: begin rgb_reg = 3'b111; end
            18'b101000101100011001: begin rgb_reg = 3'b111; end
            18'b101000101100011100: begin rgb_reg = 3'b111; end
            18'b101000101100011101: begin rgb_reg = 3'b111; end
            18'b101000101100011110: begin rgb_reg = 3'b111; end
            18'b101000101100110011: begin rgb_reg = 3'b111; end
            18'b101000101100110100: begin rgb_reg = 3'b111; end
            18'b101000101100111100: begin rgb_reg = 3'b111; end
            18'b101000101100111101: begin rgb_reg = 3'b111; end
            18'b101000110010111110: begin rgb_reg = 3'b111; end
            18'b101000110010111111: begin rgb_reg = 3'b111; end
            18'b101000110011000000: begin rgb_reg = 3'b111; end
            18'b101000110011000001: begin rgb_reg = 3'b111; end
            18'b101000110011000010: begin rgb_reg = 3'b111; end
            18'b101000110011000011: begin rgb_reg = 3'b111; end
            18'b101000110011000100: begin rgb_reg = 3'b111; end
            18'b101000110011000101: begin rgb_reg = 3'b111; end
            18'b101000110011000110: begin rgb_reg = 3'b111; end
            18'b101000110011001011: begin rgb_reg = 3'b111; end
            18'b101000110011001100: begin rgb_reg = 3'b111; end
            18'b101000110011001101: begin rgb_reg = 3'b111; end
            18'b101000110011010000: begin rgb_reg = 3'b111; end
            18'b101000110011010001: begin rgb_reg = 3'b111; end
            18'b101000110011010100: begin rgb_reg = 3'b111; end
            18'b101000110011010101: begin rgb_reg = 3'b111; end
            18'b101000110011010110: begin rgb_reg = 3'b111; end
            18'b101000110011011101: begin rgb_reg = 3'b111; end
            18'b101000110011011110: begin rgb_reg = 3'b111; end
            18'b101000110011011111: begin rgb_reg = 3'b111; end
            18'b101000110011100000: begin rgb_reg = 3'b111; end
            18'b101000110011100001: begin rgb_reg = 3'b111; end
            18'b101000110011101011: begin rgb_reg = 3'b111; end
            18'b101000110011101100: begin rgb_reg = 3'b111; end
            18'b101000110011110100: begin rgb_reg = 3'b111; end
            18'b101000110011110101: begin rgb_reg = 3'b111; end
            18'b101000110011111000: begin rgb_reg = 3'b111; end
            18'b101000110011111001: begin rgb_reg = 3'b111; end
            18'b101000110011111010: begin rgb_reg = 3'b111; end
            18'b101000110011111101: begin rgb_reg = 3'b111; end
            18'b101000110011111110: begin rgb_reg = 3'b111; end
            18'b101000110100000110: begin rgb_reg = 3'b111; end
            18'b101000110100000111: begin rgb_reg = 3'b111; end
            18'b101000110100001111: begin rgb_reg = 3'b111; end
            18'b101000110100010000: begin rgb_reg = 3'b111; end
            18'b101000110100011000: begin rgb_reg = 3'b111; end
            18'b101000110100011001: begin rgb_reg = 3'b111; end
            18'b101000110100011100: begin rgb_reg = 3'b111; end
            18'b101000110100011101: begin rgb_reg = 3'b111; end
            18'b101000110100011110: begin rgb_reg = 3'b111; end
            18'b101000110100011111: begin rgb_reg = 3'b111; end
            18'b101000110100100000: begin rgb_reg = 3'b111; end
            18'b101000110100100001: begin rgb_reg = 3'b111; end
            18'b101000110100100010: begin rgb_reg = 3'b111; end
            18'b101000110100100011: begin rgb_reg = 3'b111; end
            18'b101000110100100100: begin rgb_reg = 3'b111; end
            18'b101000110100101110: begin rgb_reg = 3'b111; end
            18'b101000110100101111: begin rgb_reg = 3'b111; end
            18'b101000110100110000: begin rgb_reg = 3'b111; end
            18'b101000110100110001: begin rgb_reg = 3'b111; end
            18'b101000110100110010: begin rgb_reg = 3'b111; end
            18'b101000110100111100: begin rgb_reg = 3'b111; end
            18'b101000110100111101: begin rgb_reg = 3'b111; end
            18'b101000111010111110: begin rgb_reg = 3'b111; end
            18'b101000111010111111: begin rgb_reg = 3'b111; end
            18'b101000111011000000: begin rgb_reg = 3'b111; end
            18'b101000111011000001: begin rgb_reg = 3'b111; end
            18'b101000111011000010: begin rgb_reg = 3'b111; end
            18'b101000111011000011: begin rgb_reg = 3'b111; end
            18'b101000111011000100: begin rgb_reg = 3'b111; end
            18'b101000111011000101: begin rgb_reg = 3'b111; end
            18'b101000111011000110: begin rgb_reg = 3'b111; end
            18'b101000111011001011: begin rgb_reg = 3'b111; end
            18'b101000111011001100: begin rgb_reg = 3'b111; end
            18'b101000111011001101: begin rgb_reg = 3'b111; end
            18'b101000111011010000: begin rgb_reg = 3'b111; end
            18'b101000111011010001: begin rgb_reg = 3'b111; end
            18'b101000111011010100: begin rgb_reg = 3'b111; end
            18'b101000111011010101: begin rgb_reg = 3'b111; end
            18'b101000111011010110: begin rgb_reg = 3'b111; end
            18'b101000111011011101: begin rgb_reg = 3'b111; end
            18'b101000111011011110: begin rgb_reg = 3'b111; end
            18'b101000111011011111: begin rgb_reg = 3'b111; end
            18'b101000111011100000: begin rgb_reg = 3'b111; end
            18'b101000111011100001: begin rgb_reg = 3'b111; end
            18'b101000111011101011: begin rgb_reg = 3'b111; end
            18'b101000111011101100: begin rgb_reg = 3'b111; end
            18'b101000111011110100: begin rgb_reg = 3'b111; end
            18'b101000111011110101: begin rgb_reg = 3'b111; end
            18'b101000111011111000: begin rgb_reg = 3'b111; end
            18'b101000111011111001: begin rgb_reg = 3'b111; end
            18'b101000111011111010: begin rgb_reg = 3'b111; end
            18'b101000111011111101: begin rgb_reg = 3'b111; end
            18'b101000111011111110: begin rgb_reg = 3'b111; end
            18'b101000111100000110: begin rgb_reg = 3'b111; end
            18'b101000111100000111: begin rgb_reg = 3'b111; end
            18'b101000111100001111: begin rgb_reg = 3'b111; end
            18'b101000111100010000: begin rgb_reg = 3'b111; end
            18'b101000111100011000: begin rgb_reg = 3'b111; end
            18'b101000111100011001: begin rgb_reg = 3'b111; end
            18'b101000111100011100: begin rgb_reg = 3'b111; end
            18'b101000111100011101: begin rgb_reg = 3'b111; end
            18'b101000111100011110: begin rgb_reg = 3'b111; end
            18'b101000111100011111: begin rgb_reg = 3'b111; end
            18'b101000111100100000: begin rgb_reg = 3'b111; end
            18'b101000111100100001: begin rgb_reg = 3'b111; end
            18'b101000111100100010: begin rgb_reg = 3'b111; end
            18'b101000111100100011: begin rgb_reg = 3'b111; end
            18'b101000111100100100: begin rgb_reg = 3'b111; end
            18'b101000111100101110: begin rgb_reg = 3'b111; end
            18'b101000111100101111: begin rgb_reg = 3'b111; end
            18'b101000111100110000: begin rgb_reg = 3'b111; end
            18'b101000111100110001: begin rgb_reg = 3'b111; end
            18'b101000111100110010: begin rgb_reg = 3'b111; end
            18'b101000111100111100: begin rgb_reg = 3'b111; end
            18'b101000111100111101: begin rgb_reg = 3'b111; end
            18'b101001000010111110: begin rgb_reg = 3'b111; end
            18'b101001000010111111: begin rgb_reg = 3'b111; end
            18'b101001000011000111: begin rgb_reg = 3'b111; end
            18'b101001000011001000: begin rgb_reg = 3'b111; end
            18'b101001000011001011: begin rgb_reg = 3'b111; end
            18'b101001000011001100: begin rgb_reg = 3'b111; end
            18'b101001000011001101: begin rgb_reg = 3'b111; end
            18'b101001000011001110: begin rgb_reg = 3'b111; end
            18'b101001000011001111: begin rgb_reg = 3'b111; end
            18'b101001000011010100: begin rgb_reg = 3'b111; end
            18'b101001000011010101: begin rgb_reg = 3'b111; end
            18'b101001000011010110: begin rgb_reg = 3'b111; end
            18'b101001000011100010: begin rgb_reg = 3'b111; end
            18'b101001000011100011: begin rgb_reg = 3'b111; end
            18'b101001000011101011: begin rgb_reg = 3'b111; end
            18'b101001000011101100: begin rgb_reg = 3'b111; end
            18'b101001000011110100: begin rgb_reg = 3'b111; end
            18'b101001000011110101: begin rgb_reg = 3'b111; end
            18'b101001000011110110: begin rgb_reg = 3'b111; end
            18'b101001000011110111: begin rgb_reg = 3'b111; end
            18'b101001000011111101: begin rgb_reg = 3'b111; end
            18'b101001000011111110: begin rgb_reg = 3'b111; end
            18'b101001000100000110: begin rgb_reg = 3'b111; end
            18'b101001000100000111: begin rgb_reg = 3'b111; end
            18'b101001000100001111: begin rgb_reg = 3'b111; end
            18'b101001000100010000: begin rgb_reg = 3'b111; end
            18'b101001000100010001: begin rgb_reg = 3'b111; end
            18'b101001000100010010: begin rgb_reg = 3'b111; end
            18'b101001000100010011: begin rgb_reg = 3'b111; end
            18'b101001000100010100: begin rgb_reg = 3'b111; end
            18'b101001000100010101: begin rgb_reg = 3'b111; end
            18'b101001000100010110: begin rgb_reg = 3'b111; end
            18'b101001000100010111: begin rgb_reg = 3'b111; end
            18'b101001000100011000: begin rgb_reg = 3'b111; end
            18'b101001000100011001: begin rgb_reg = 3'b111; end
            18'b101001000100011100: begin rgb_reg = 3'b111; end
            18'b101001000100011101: begin rgb_reg = 3'b111; end
            18'b101001000100011110: begin rgb_reg = 3'b111; end
            18'b101001000100100101: begin rgb_reg = 3'b111; end
            18'b101001000100100110: begin rgb_reg = 3'b111; end
            18'b101001000100100111: begin rgb_reg = 3'b111; end
            18'b101001000100101100: begin rgb_reg = 3'b111; end
            18'b101001000100101101: begin rgb_reg = 3'b111; end
            18'b101001000100111100: begin rgb_reg = 3'b111; end
            18'b101001000100111101: begin rgb_reg = 3'b111; end
            18'b101001001010111110: begin rgb_reg = 3'b111; end
            18'b101001001010111111: begin rgb_reg = 3'b111; end
            18'b101001001011000111: begin rgb_reg = 3'b111; end
            18'b101001001011001000: begin rgb_reg = 3'b111; end
            18'b101001001011001011: begin rgb_reg = 3'b111; end
            18'b101001001011001100: begin rgb_reg = 3'b111; end
            18'b101001001011001101: begin rgb_reg = 3'b111; end
            18'b101001001011001110: begin rgb_reg = 3'b111; end
            18'b101001001011001111: begin rgb_reg = 3'b111; end
            18'b101001001011010100: begin rgb_reg = 3'b111; end
            18'b101001001011010101: begin rgb_reg = 3'b111; end
            18'b101001001011010110: begin rgb_reg = 3'b111; end
            18'b101001001011100010: begin rgb_reg = 3'b111; end
            18'b101001001011100011: begin rgb_reg = 3'b111; end
            18'b101001001011101011: begin rgb_reg = 3'b111; end
            18'b101001001011101100: begin rgb_reg = 3'b111; end
            18'b101001001011110100: begin rgb_reg = 3'b111; end
            18'b101001001011110101: begin rgb_reg = 3'b111; end
            18'b101001001011110110: begin rgb_reg = 3'b111; end
            18'b101001001011110111: begin rgb_reg = 3'b111; end
            18'b101001001011111101: begin rgb_reg = 3'b111; end
            18'b101001001011111110: begin rgb_reg = 3'b111; end
            18'b101001001100000110: begin rgb_reg = 3'b111; end
            18'b101001001100000111: begin rgb_reg = 3'b111; end
            18'b101001001100001111: begin rgb_reg = 3'b111; end
            18'b101001001100010000: begin rgb_reg = 3'b111; end
            18'b101001001100010001: begin rgb_reg = 3'b111; end
            18'b101001001100010010: begin rgb_reg = 3'b111; end
            18'b101001001100010011: begin rgb_reg = 3'b111; end
            18'b101001001100010100: begin rgb_reg = 3'b111; end
            18'b101001001100010101: begin rgb_reg = 3'b111; end
            18'b101001001100010110: begin rgb_reg = 3'b111; end
            18'b101001001100010111: begin rgb_reg = 3'b111; end
            18'b101001001100011000: begin rgb_reg = 3'b111; end
            18'b101001001100011001: begin rgb_reg = 3'b111; end
            18'b101001001100011100: begin rgb_reg = 3'b111; end
            18'b101001001100011101: begin rgb_reg = 3'b111; end
            18'b101001001100011110: begin rgb_reg = 3'b111; end
            18'b101001001100100101: begin rgb_reg = 3'b111; end
            18'b101001001100100110: begin rgb_reg = 3'b111; end
            18'b101001001100100111: begin rgb_reg = 3'b111; end
            18'b101001001100101100: begin rgb_reg = 3'b111; end
            18'b101001001100101101: begin rgb_reg = 3'b111; end
            18'b101001001100111100: begin rgb_reg = 3'b111; end
            18'b101001001100111101: begin rgb_reg = 3'b111; end
            18'b101001010010111110: begin rgb_reg = 3'b111; end
            18'b101001010010111111: begin rgb_reg = 3'b111; end
            18'b101001010011000111: begin rgb_reg = 3'b111; end
            18'b101001010011001000: begin rgb_reg = 3'b111; end
            18'b101001010011001011: begin rgb_reg = 3'b111; end
            18'b101001010011001100: begin rgb_reg = 3'b111; end
            18'b101001010011001101: begin rgb_reg = 3'b111; end
            18'b101001010011010100: begin rgb_reg = 3'b111; end
            18'b101001010011010101: begin rgb_reg = 3'b111; end
            18'b101001010011010110: begin rgb_reg = 3'b111; end
            18'b101001010011011001: begin rgb_reg = 3'b111; end
            18'b101001010011011010: begin rgb_reg = 3'b111; end
            18'b101001010011100010: begin rgb_reg = 3'b111; end
            18'b101001010011100011: begin rgb_reg = 3'b111; end
            18'b101001010011101011: begin rgb_reg = 3'b111; end
            18'b101001010011101100: begin rgb_reg = 3'b111; end
            18'b101001010011110100: begin rgb_reg = 3'b111; end
            18'b101001010011110101: begin rgb_reg = 3'b111; end
            18'b101001010011111101: begin rgb_reg = 3'b111; end
            18'b101001010011111110: begin rgb_reg = 3'b111; end
            18'b101001010100000110: begin rgb_reg = 3'b111; end
            18'b101001010100000111: begin rgb_reg = 3'b111; end
            18'b101001010100010111: begin rgb_reg = 3'b111; end
            18'b101001010100011000: begin rgb_reg = 3'b111; end
            18'b101001010100011001: begin rgb_reg = 3'b111; end
            18'b101001010100011100: begin rgb_reg = 3'b111; end
            18'b101001010100011101: begin rgb_reg = 3'b111; end
            18'b101001010100011110: begin rgb_reg = 3'b111; end
            18'b101001010100100101: begin rgb_reg = 3'b111; end
            18'b101001010100100110: begin rgb_reg = 3'b111; end
            18'b101001010100100111: begin rgb_reg = 3'b111; end
            18'b101001010100101010: begin rgb_reg = 3'b111; end
            18'b101001010100101011: begin rgb_reg = 3'b111; end
            18'b101001010100111100: begin rgb_reg = 3'b111; end
            18'b101001010100111101: begin rgb_reg = 3'b111; end
            18'b101001011010111110: begin rgb_reg = 3'b111; end
            18'b101001011010111111: begin rgb_reg = 3'b111; end
            18'b101001011011000111: begin rgb_reg = 3'b111; end
            18'b101001011011001000: begin rgb_reg = 3'b111; end
            18'b101001011011001011: begin rgb_reg = 3'b111; end
            18'b101001011011001100: begin rgb_reg = 3'b111; end
            18'b101001011011001101: begin rgb_reg = 3'b111; end
            18'b101001011011010100: begin rgb_reg = 3'b111; end
            18'b101001011011010101: begin rgb_reg = 3'b111; end
            18'b101001011011010110: begin rgb_reg = 3'b111; end
            18'b101001011011011001: begin rgb_reg = 3'b111; end
            18'b101001011011011010: begin rgb_reg = 3'b111; end
            18'b101001011011100010: begin rgb_reg = 3'b111; end
            18'b101001011011100011: begin rgb_reg = 3'b111; end
            18'b101001011011101011: begin rgb_reg = 3'b111; end
            18'b101001011011101100: begin rgb_reg = 3'b111; end
            18'b101001011011110100: begin rgb_reg = 3'b111; end
            18'b101001011011110101: begin rgb_reg = 3'b111; end
            18'b101001011011111101: begin rgb_reg = 3'b111; end
            18'b101001011011111110: begin rgb_reg = 3'b111; end
            18'b101001011100000110: begin rgb_reg = 3'b111; end
            18'b101001011100000111: begin rgb_reg = 3'b111; end
            18'b101001011100011000: begin rgb_reg = 3'b111; end
            18'b101001011100011001: begin rgb_reg = 3'b111; end
            18'b101001011100011100: begin rgb_reg = 3'b111; end
            18'b101001011100011101: begin rgb_reg = 3'b111; end
            18'b101001011100011110: begin rgb_reg = 3'b111; end
            18'b101001011100100101: begin rgb_reg = 3'b111; end
            18'b101001011100100110: begin rgb_reg = 3'b111; end
            18'b101001011100100111: begin rgb_reg = 3'b111; end
            18'b101001011100101010: begin rgb_reg = 3'b111; end
            18'b101001011100101011: begin rgb_reg = 3'b111; end
            18'b101001011100111100: begin rgb_reg = 3'b111; end
            18'b101001011100111101: begin rgb_reg = 3'b111; end
            18'b101001100010111110: begin rgb_reg = 3'b111; end
            18'b101001100010111111: begin rgb_reg = 3'b111; end
            18'b101001100011000000: begin rgb_reg = 3'b111; end
            18'b101001100011000001: begin rgb_reg = 3'b111; end
            18'b101001100011000010: begin rgb_reg = 3'b111; end
            18'b101001100011000011: begin rgb_reg = 3'b111; end
            18'b101001100011000100: begin rgb_reg = 3'b111; end
            18'b101001100011000101: begin rgb_reg = 3'b111; end
            18'b101001100011000110: begin rgb_reg = 3'b111; end
            18'b101001100011000111: begin rgb_reg = 3'b111; end
            18'b101001100011001000: begin rgb_reg = 3'b111; end
            18'b101001100011001100: begin rgb_reg = 3'b111; end
            18'b101001100011001101: begin rgb_reg = 3'b111; end
            18'b101001100011001110: begin rgb_reg = 3'b111; end
            18'b101001100011001111: begin rgb_reg = 3'b111; end
            18'b101001100011010000: begin rgb_reg = 3'b111; end
            18'b101001100011010001: begin rgb_reg = 3'b111; end
            18'b101001100011010010: begin rgb_reg = 3'b111; end
            18'b101001100011010011: begin rgb_reg = 3'b111; end
            18'b101001100011010100: begin rgb_reg = 3'b111; end
            18'b101001100011010101: begin rgb_reg = 3'b111; end
            18'b101001100011011001: begin rgb_reg = 3'b111; end
            18'b101001100011011010: begin rgb_reg = 3'b111; end
            18'b101001100011011011: begin rgb_reg = 3'b111; end
            18'b101001100011011100: begin rgb_reg = 3'b111; end
            18'b101001100011011101: begin rgb_reg = 3'b111; end
            18'b101001100011011110: begin rgb_reg = 3'b111; end
            18'b101001100011011111: begin rgb_reg = 3'b111; end
            18'b101001100011100000: begin rgb_reg = 3'b111; end
            18'b101001100011100001: begin rgb_reg = 3'b111; end
            18'b101001100011100010: begin rgb_reg = 3'b111; end
            18'b101001100011100011: begin rgb_reg = 3'b111; end
            18'b101001100011100111: begin rgb_reg = 3'b111; end
            18'b101001100011101000: begin rgb_reg = 3'b111; end
            18'b101001100011101001: begin rgb_reg = 3'b111; end
            18'b101001100011101010: begin rgb_reg = 3'b111; end
            18'b101001100011101011: begin rgb_reg = 3'b111; end
            18'b101001100011101100: begin rgb_reg = 3'b111; end
            18'b101001100011101101: begin rgb_reg = 3'b111; end
            18'b101001100011101110: begin rgb_reg = 3'b111; end
            18'b101001100011101111: begin rgb_reg = 3'b111; end
            18'b101001100011110000: begin rgb_reg = 3'b111; end
            18'b101001100011110100: begin rgb_reg = 3'b111; end
            18'b101001100011110101: begin rgb_reg = 3'b111; end
            18'b101001100011110110: begin rgb_reg = 3'b111; end
            18'b101001100011110111: begin rgb_reg = 3'b111; end
            18'b101001100011111000: begin rgb_reg = 3'b111; end
            18'b101001100011111001: begin rgb_reg = 3'b111; end
            18'b101001100011111010: begin rgb_reg = 3'b111; end
            18'b101001100011111011: begin rgb_reg = 3'b111; end
            18'b101001100011111100: begin rgb_reg = 3'b111; end
            18'b101001100011111101: begin rgb_reg = 3'b111; end
            18'b101001100011111110: begin rgb_reg = 3'b111; end
            18'b101001100100000010: begin rgb_reg = 3'b111; end
            18'b101001100100000011: begin rgb_reg = 3'b111; end
            18'b101001100100000100: begin rgb_reg = 3'b111; end
            18'b101001100100000101: begin rgb_reg = 3'b111; end
            18'b101001100100000110: begin rgb_reg = 3'b111; end
            18'b101001100100000111: begin rgb_reg = 3'b111; end
            18'b101001100100001000: begin rgb_reg = 3'b111; end
            18'b101001100100001001: begin rgb_reg = 3'b111; end
            18'b101001100100001010: begin rgb_reg = 3'b111; end
            18'b101001100100001011: begin rgb_reg = 3'b111; end
            18'b101001100100011000: begin rgb_reg = 3'b111; end
            18'b101001100100011001: begin rgb_reg = 3'b111; end
            18'b101001100100011101: begin rgb_reg = 3'b111; end
            18'b101001100100011110: begin rgb_reg = 3'b111; end
            18'b101001100100011111: begin rgb_reg = 3'b111; end
            18'b101001100100100000: begin rgb_reg = 3'b111; end
            18'b101001100100100001: begin rgb_reg = 3'b111; end
            18'b101001100100100010: begin rgb_reg = 3'b111; end
            18'b101001100100100011: begin rgb_reg = 3'b111; end
            18'b101001100100100100: begin rgb_reg = 3'b111; end
            18'b101001100100100101: begin rgb_reg = 3'b111; end
            18'b101001100100100110: begin rgb_reg = 3'b111; end
            18'b101001100100101010: begin rgb_reg = 3'b111; end
            18'b101001100100101011: begin rgb_reg = 3'b111; end
            18'b101001100100101100: begin rgb_reg = 3'b111; end
            18'b101001100100101101: begin rgb_reg = 3'b111; end
            18'b101001100100101110: begin rgb_reg = 3'b111; end
            18'b101001100100101111: begin rgb_reg = 3'b111; end
            18'b101001100100110000: begin rgb_reg = 3'b111; end
            18'b101001100100110001: begin rgb_reg = 3'b111; end
            18'b101001100100110010: begin rgb_reg = 3'b111; end
            18'b101001100100110011: begin rgb_reg = 3'b111; end
            18'b101001100100110100: begin rgb_reg = 3'b111; end
            18'b101001100100111000: begin rgb_reg = 3'b111; end
            18'b101001100100111001: begin rgb_reg = 3'b111; end
            18'b101001100100111010: begin rgb_reg = 3'b111; end
            18'b101001100100111011: begin rgb_reg = 3'b111; end
            18'b101001100100111100: begin rgb_reg = 3'b111; end
            18'b101001100100111101: begin rgb_reg = 3'b111; end
            18'b101001100100111110: begin rgb_reg = 3'b111; end
            18'b101001100100111111: begin rgb_reg = 3'b111; end
            18'b101001100101000000: begin rgb_reg = 3'b111; end
            18'b101001100101000001: begin rgb_reg = 3'b111; end
            18'b101001101011000000: begin rgb_reg = 3'b111; end
            18'b101001101011000001: begin rgb_reg = 3'b111; end
            18'b101001101011000010: begin rgb_reg = 3'b111; end
            18'b101001101011000011: begin rgb_reg = 3'b111; end
            18'b101001101011000100: begin rgb_reg = 3'b111; end
            18'b101001101011000101: begin rgb_reg = 3'b111; end
            18'b101001101011000110: begin rgb_reg = 3'b111; end
            18'b101001101011001101: begin rgb_reg = 3'b111; end
            18'b101001101011001110: begin rgb_reg = 3'b111; end
            18'b101001101011001111: begin rgb_reg = 3'b111; end
            18'b101001101011010000: begin rgb_reg = 3'b111; end
            18'b101001101011010001: begin rgb_reg = 3'b111; end
            18'b101001101011010010: begin rgb_reg = 3'b111; end
            18'b101001101011010011: begin rgb_reg = 3'b111; end
            18'b101001101011011011: begin rgb_reg = 3'b111; end
            18'b101001101011011100: begin rgb_reg = 3'b111; end
            18'b101001101011011101: begin rgb_reg = 3'b111; end
            18'b101001101011011110: begin rgb_reg = 3'b111; end
            18'b101001101011011111: begin rgb_reg = 3'b111; end
            18'b101001101011100000: begin rgb_reg = 3'b111; end
            18'b101001101011100001: begin rgb_reg = 3'b111; end
            18'b101001101011100110: begin rgb_reg = 3'b111; end
            18'b101001101011100111: begin rgb_reg = 3'b111; end
            18'b101001101011101000: begin rgb_reg = 3'b111; end
            18'b101001101011101001: begin rgb_reg = 3'b111; end
            18'b101001101011101010: begin rgb_reg = 3'b111; end
            18'b101001101011101011: begin rgb_reg = 3'b111; end
            18'b101001101011101100: begin rgb_reg = 3'b111; end
            18'b101001101011101101: begin rgb_reg = 3'b111; end
            18'b101001101011101110: begin rgb_reg = 3'b111; end
            18'b101001101011101111: begin rgb_reg = 3'b111; end
            18'b101001101011110000: begin rgb_reg = 3'b111; end
            18'b101001101011110001: begin rgb_reg = 3'b111; end
            18'b101001101011110110: begin rgb_reg = 3'b111; end
            18'b101001101011110111: begin rgb_reg = 3'b111; end
            18'b101001101011111000: begin rgb_reg = 3'b111; end
            18'b101001101011111001: begin rgb_reg = 3'b111; end
            18'b101001101011111010: begin rgb_reg = 3'b111; end
            18'b101001101011111011: begin rgb_reg = 3'b111; end
            18'b101001101011111100: begin rgb_reg = 3'b111; end
            18'b101001101100000001: begin rgb_reg = 3'b111; end
            18'b101001101100000010: begin rgb_reg = 3'b111; end
            18'b101001101100000011: begin rgb_reg = 3'b111; end
            18'b101001101100000100: begin rgb_reg = 3'b111; end
            18'b101001101100000101: begin rgb_reg = 3'b111; end
            18'b101001101100000110: begin rgb_reg = 3'b111; end
            18'b101001101100000111: begin rgb_reg = 3'b111; end
            18'b101001101100001000: begin rgb_reg = 3'b111; end
            18'b101001101100001001: begin rgb_reg = 3'b111; end
            18'b101001101100001010: begin rgb_reg = 3'b111; end
            18'b101001101100001011: begin rgb_reg = 3'b111; end
            18'b101001101100001100: begin rgb_reg = 3'b111; end
            18'b101001101100011000: begin rgb_reg = 3'b111; end
            18'b101001101100011001: begin rgb_reg = 3'b111; end
            18'b101001101100011110: begin rgb_reg = 3'b111; end
            18'b101001101100011111: begin rgb_reg = 3'b111; end
            18'b101001101100100000: begin rgb_reg = 3'b111; end
            18'b101001101100100001: begin rgb_reg = 3'b111; end
            18'b101001101100100010: begin rgb_reg = 3'b111; end
            18'b101001101100100011: begin rgb_reg = 3'b111; end
            18'b101001101100100100: begin rgb_reg = 3'b111; end
            18'b101001101100101010: begin rgb_reg = 3'b111; end
            18'b101001101100101011: begin rgb_reg = 3'b111; end
            18'b101001101100101100: begin rgb_reg = 3'b111; end
            18'b101001101100101101: begin rgb_reg = 3'b111; end
            18'b101001101100101110: begin rgb_reg = 3'b111; end
            18'b101001101100101111: begin rgb_reg = 3'b111; end
            18'b101001101100110000: begin rgb_reg = 3'b111; end
            18'b101001101100110001: begin rgb_reg = 3'b111; end
            18'b101001101100110010: begin rgb_reg = 3'b111; end
            18'b101001101100110011: begin rgb_reg = 3'b111; end
            18'b101001101100110100: begin rgb_reg = 3'b111; end
            18'b101001101100110111: begin rgb_reg = 3'b111; end
            18'b101001101100111000: begin rgb_reg = 3'b111; end
            18'b101001101100111001: begin rgb_reg = 3'b111; end
            18'b101001101100111010: begin rgb_reg = 3'b111; end
            18'b101001101100111011: begin rgb_reg = 3'b111; end
            18'b101001101100111100: begin rgb_reg = 3'b111; end
            18'b101001101100111101: begin rgb_reg = 3'b111; end
            18'b101001101100111110: begin rgb_reg = 3'b111; end
            18'b101001101100111111: begin rgb_reg = 3'b111; end
            18'b101001101101000000: begin rgb_reg = 3'b111; end
            18'b101001101101000001: begin rgb_reg = 3'b111; end
            18'b101001101101000010: begin rgb_reg = 3'b111; end
            18'b101001110011000000: begin rgb_reg = 3'b111; end
            18'b101001110011000001: begin rgb_reg = 3'b111; end
            18'b101001110011000010: begin rgb_reg = 3'b111; end
            18'b101001110011000011: begin rgb_reg = 3'b111; end
            18'b101001110011000100: begin rgb_reg = 3'b111; end
            18'b101001110011000101: begin rgb_reg = 3'b111; end
            18'b101001110011000110: begin rgb_reg = 3'b111; end
            18'b101001110011001110: begin rgb_reg = 3'b111; end
            18'b101001110011001111: begin rgb_reg = 3'b111; end
            18'b101001110011010000: begin rgb_reg = 3'b111; end
            18'b101001110011010001: begin rgb_reg = 3'b111; end
            18'b101001110011010010: begin rgb_reg = 3'b111; end
            18'b101001110011010011: begin rgb_reg = 3'b111; end
            18'b101001110011011011: begin rgb_reg = 3'b111; end
            18'b101001110011011100: begin rgb_reg = 3'b111; end
            18'b101001110011011101: begin rgb_reg = 3'b111; end
            18'b101001110011011110: begin rgb_reg = 3'b111; end
            18'b101001110011011111: begin rgb_reg = 3'b111; end
            18'b101001110011100000: begin rgb_reg = 3'b111; end
            18'b101001110011100001: begin rgb_reg = 3'b111; end
            18'b101001110011100110: begin rgb_reg = 3'b111; end
            18'b101001110011100111: begin rgb_reg = 3'b111; end
            18'b101001110011101000: begin rgb_reg = 3'b111; end
            18'b101001110011101001: begin rgb_reg = 3'b111; end
            18'b101001110011101010: begin rgb_reg = 3'b111; end
            18'b101001110011101011: begin rgb_reg = 3'b111; end
            18'b101001110011101100: begin rgb_reg = 3'b111; end
            18'b101001110011101101: begin rgb_reg = 3'b111; end
            18'b101001110011101110: begin rgb_reg = 3'b111; end
            18'b101001110011101111: begin rgb_reg = 3'b111; end
            18'b101001110011110000: begin rgb_reg = 3'b111; end
            18'b101001110011110110: begin rgb_reg = 3'b111; end
            18'b101001110011110111: begin rgb_reg = 3'b111; end
            18'b101001110011111000: begin rgb_reg = 3'b111; end
            18'b101001110011111001: begin rgb_reg = 3'b111; end
            18'b101001110011111010: begin rgb_reg = 3'b111; end
            18'b101001110011111011: begin rgb_reg = 3'b111; end
            18'b101001110011111100: begin rgb_reg = 3'b111; end
            18'b101001110100000001: begin rgb_reg = 3'b111; end
            18'b101001110100000010: begin rgb_reg = 3'b111; end
            18'b101001110100000011: begin rgb_reg = 3'b111; end
            18'b101001110100000100: begin rgb_reg = 3'b111; end
            18'b101001110100000101: begin rgb_reg = 3'b111; end
            18'b101001110100000110: begin rgb_reg = 3'b111; end
            18'b101001110100000111: begin rgb_reg = 3'b111; end
            18'b101001110100001000: begin rgb_reg = 3'b111; end
            18'b101001110100001001: begin rgb_reg = 3'b111; end
            18'b101001110100001010: begin rgb_reg = 3'b111; end
            18'b101001110100001011: begin rgb_reg = 3'b111; end
            18'b101001110100011000: begin rgb_reg = 3'b111; end
            18'b101001110100011001: begin rgb_reg = 3'b111; end
            18'b101001110100011111: begin rgb_reg = 3'b111; end
            18'b101001110100100000: begin rgb_reg = 3'b111; end
            18'b101001110100100001: begin rgb_reg = 3'b111; end
            18'b101001110100100010: begin rgb_reg = 3'b111; end
            18'b101001110100100011: begin rgb_reg = 3'b111; end
            18'b101001110100100100: begin rgb_reg = 3'b111; end
            18'b101001110100101010: begin rgb_reg = 3'b111; end
            18'b101001110100101011: begin rgb_reg = 3'b111; end
            18'b101001110100101100: begin rgb_reg = 3'b111; end
            18'b101001110100101101: begin rgb_reg = 3'b111; end
            18'b101001110100101110: begin rgb_reg = 3'b111; end
            18'b101001110100101111: begin rgb_reg = 3'b111; end
            18'b101001110100110000: begin rgb_reg = 3'b111; end
            18'b101001110100110001: begin rgb_reg = 3'b111; end
            18'b101001110100110010: begin rgb_reg = 3'b111; end
            18'b101001110100110011: begin rgb_reg = 3'b111; end
            18'b101001110100110100: begin rgb_reg = 3'b111; end
            18'b101001110100110111: begin rgb_reg = 3'b111; end
            18'b101001110100111000: begin rgb_reg = 3'b111; end
            18'b101001110100111001: begin rgb_reg = 3'b111; end
            18'b101001110100111010: begin rgb_reg = 3'b111; end
            18'b101001110100111011: begin rgb_reg = 3'b111; end
            18'b101001110100111100: begin rgb_reg = 3'b111; end
            18'b101001110100111101: begin rgb_reg = 3'b111; end
            18'b101001110100111110: begin rgb_reg = 3'b111; end
            18'b101001110100111111: begin rgb_reg = 3'b111; end
            18'b101001110101000000: begin rgb_reg = 3'b111; end
            18'b101001110101000001: begin rgb_reg = 3'b111; end
            18'b101010101010001001: begin rgb_reg = 3'b111; end
            18'b101010101010001010: begin rgb_reg = 3'b111; end
            18'b101010101010010001: begin rgb_reg = 3'b111; end
            18'b101010101010010010: begin rgb_reg = 3'b111; end
            18'b101010101010100011: begin rgb_reg = 3'b111; end
            18'b101010101010100100: begin rgb_reg = 3'b111; end
            18'b101010101010101001: begin rgb_reg = 3'b111; end
            18'b101010101010101010: begin rgb_reg = 3'b111; end
            18'b101010101011001101: begin rgb_reg = 3'b111; end
            18'b101010101011001110: begin rgb_reg = 3'b111; end
            18'b101010101011111101: begin rgb_reg = 3'b111; end
            18'b101010101011111110: begin rgb_reg = 3'b111; end
            18'b101010101100000101: begin rgb_reg = 3'b111; end
            18'b101010101100000110: begin rgb_reg = 3'b111; end
            18'b101010101100001001: begin rgb_reg = 3'b111; end
            18'b101010101100001010: begin rgb_reg = 3'b111; end
            18'b101010101101001011: begin rgb_reg = 3'b111; end
            18'b101010101101001100: begin rgb_reg = 3'b111; end
            18'b101010101101010001: begin rgb_reg = 3'b111; end
            18'b101010101101010010: begin rgb_reg = 3'b111; end
            18'b101010101101011101: begin rgb_reg = 3'b111; end
            18'b101010101101011110: begin rgb_reg = 3'b111; end
            18'b101010110010001001: begin rgb_reg = 3'b111; end
            18'b101010110010001010: begin rgb_reg = 3'b111; end
            18'b101010110010010001: begin rgb_reg = 3'b111; end
            18'b101010110010010010: begin rgb_reg = 3'b111; end
            18'b101010110010100011: begin rgb_reg = 3'b111; end
            18'b101010110010100100: begin rgb_reg = 3'b111; end
            18'b101010110010101001: begin rgb_reg = 3'b111; end
            18'b101010110010101010: begin rgb_reg = 3'b111; end
            18'b101010110011001101: begin rgb_reg = 3'b111; end
            18'b101010110011001110: begin rgb_reg = 3'b111; end
            18'b101010110011111101: begin rgb_reg = 3'b111; end
            18'b101010110011111110: begin rgb_reg = 3'b111; end
            18'b101010110100000101: begin rgb_reg = 3'b111; end
            18'b101010110100000110: begin rgb_reg = 3'b111; end
            18'b101010110100001001: begin rgb_reg = 3'b111; end
            18'b101010110100001010: begin rgb_reg = 3'b111; end
            18'b101010110101001011: begin rgb_reg = 3'b111; end
            18'b101010110101001100: begin rgb_reg = 3'b111; end
            18'b101010110101010001: begin rgb_reg = 3'b111; end
            18'b101010110101010010: begin rgb_reg = 3'b111; end
            18'b101010110101011101: begin rgb_reg = 3'b111; end
            18'b101010110101011110: begin rgb_reg = 3'b111; end
            18'b101010111010001001: begin rgb_reg = 3'b111; end
            18'b101010111010001010: begin rgb_reg = 3'b111; end
            18'b101010111010001011: begin rgb_reg = 3'b111; end
            18'b101010111010001100: begin rgb_reg = 3'b111; end
            18'b101010111010010001: begin rgb_reg = 3'b111; end
            18'b101010111010010010: begin rgb_reg = 3'b111; end
            18'b101010111010100001: begin rgb_reg = 3'b111; end
            18'b101010111010100010: begin rgb_reg = 3'b111; end
            18'b101010111010100011: begin rgb_reg = 3'b111; end
            18'b101010111010100100: begin rgb_reg = 3'b111; end
            18'b101010111010100101: begin rgb_reg = 3'b111; end
            18'b101010111010100110: begin rgb_reg = 3'b111; end
            18'b101010111010101001: begin rgb_reg = 3'b111; end
            18'b101010111010101010: begin rgb_reg = 3'b111; end
            18'b101010111011001101: begin rgb_reg = 3'b111; end
            18'b101010111011001110: begin rgb_reg = 3'b111; end
            18'b101010111011111101: begin rgb_reg = 3'b111; end
            18'b101010111011111110: begin rgb_reg = 3'b111; end
            18'b101010111011111111: begin rgb_reg = 3'b111; end
            18'b101010111100000000: begin rgb_reg = 3'b111; end
            18'b101010111100000101: begin rgb_reg = 3'b111; end
            18'b101010111100000110: begin rgb_reg = 3'b111; end
            18'b101010111101001001: begin rgb_reg = 3'b111; end
            18'b101010111101001010: begin rgb_reg = 3'b111; end
            18'b101010111101001011: begin rgb_reg = 3'b111; end
            18'b101010111101001100: begin rgb_reg = 3'b111; end
            18'b101010111101001101: begin rgb_reg = 3'b111; end
            18'b101010111101001110: begin rgb_reg = 3'b111; end
            18'b101010111101010001: begin rgb_reg = 3'b111; end
            18'b101010111101010010: begin rgb_reg = 3'b111; end
            18'b101011000010001001: begin rgb_reg = 3'b111; end
            18'b101011000010001010: begin rgb_reg = 3'b111; end
            18'b101011000010001011: begin rgb_reg = 3'b111; end
            18'b101011000010001100: begin rgb_reg = 3'b111; end
            18'b101011000010010001: begin rgb_reg = 3'b111; end
            18'b101011000010010010: begin rgb_reg = 3'b111; end
            18'b101011000010100001: begin rgb_reg = 3'b111; end
            18'b101011000010100010: begin rgb_reg = 3'b111; end
            18'b101011000010100011: begin rgb_reg = 3'b111; end
            18'b101011000010100100: begin rgb_reg = 3'b111; end
            18'b101011000010100101: begin rgb_reg = 3'b111; end
            18'b101011000010100110: begin rgb_reg = 3'b111; end
            18'b101011000010101001: begin rgb_reg = 3'b111; end
            18'b101011000010101010: begin rgb_reg = 3'b111; end
            18'b101011000011001101: begin rgb_reg = 3'b111; end
            18'b101011000011001110: begin rgb_reg = 3'b111; end
            18'b101011000011111101: begin rgb_reg = 3'b111; end
            18'b101011000011111110: begin rgb_reg = 3'b111; end
            18'b101011000011111111: begin rgb_reg = 3'b111; end
            18'b101011000100000000: begin rgb_reg = 3'b111; end
            18'b101011000100000101: begin rgb_reg = 3'b111; end
            18'b101011000100000110: begin rgb_reg = 3'b111; end
            18'b101011000101001001: begin rgb_reg = 3'b111; end
            18'b101011000101001010: begin rgb_reg = 3'b111; end
            18'b101011000101001011: begin rgb_reg = 3'b111; end
            18'b101011000101001100: begin rgb_reg = 3'b111; end
            18'b101011000101001101: begin rgb_reg = 3'b111; end
            18'b101011000101001110: begin rgb_reg = 3'b111; end
            18'b101011000101010001: begin rgb_reg = 3'b111; end
            18'b101011000101010010: begin rgb_reg = 3'b111; end
            18'b101011001010001001: begin rgb_reg = 3'b111; end
            18'b101011001010001010: begin rgb_reg = 3'b111; end
            18'b101011001010001101: begin rgb_reg = 3'b111; end
            18'b101011001010001110: begin rgb_reg = 3'b111; end
            18'b101011001010010001: begin rgb_reg = 3'b111; end
            18'b101011001010010010: begin rgb_reg = 3'b111; end
            18'b101011001010010111: begin rgb_reg = 3'b111; end
            18'b101011001010011000: begin rgb_reg = 3'b111; end
            18'b101011001010011001: begin rgb_reg = 3'b111; end
            18'b101011001010011010: begin rgb_reg = 3'b111; end
            18'b101011001010011011: begin rgb_reg = 3'b111; end
            18'b101011001010011100: begin rgb_reg = 3'b111; end
            18'b101011001010100011: begin rgb_reg = 3'b111; end
            18'b101011001010100100: begin rgb_reg = 3'b111; end
            18'b101011001010101001: begin rgb_reg = 3'b111; end
            18'b101011001010101010: begin rgb_reg = 3'b111; end
            18'b101011001010101101: begin rgb_reg = 3'b111; end
            18'b101011001010101110: begin rgb_reg = 3'b111; end
            18'b101011001010101111: begin rgb_reg = 3'b111; end
            18'b101011001010110000: begin rgb_reg = 3'b111; end
            18'b101011001010110111: begin rgb_reg = 3'b111; end
            18'b101011001010111000: begin rgb_reg = 3'b111; end
            18'b101011001010111001: begin rgb_reg = 3'b111; end
            18'b101011001010111010: begin rgb_reg = 3'b111; end
            18'b101011001010111011: begin rgb_reg = 3'b111; end
            18'b101011001010111100: begin rgb_reg = 3'b111; end
            18'b101011001011000001: begin rgb_reg = 3'b111; end
            18'b101011001011000010: begin rgb_reg = 3'b111; end
            18'b101011001011000101: begin rgb_reg = 3'b111; end
            18'b101011001011000110: begin rgb_reg = 3'b111; end
            18'b101011001011000111: begin rgb_reg = 3'b111; end
            18'b101011001011001000: begin rgb_reg = 3'b111; end
            18'b101011001011001101: begin rgb_reg = 3'b111; end
            18'b101011001011001110: begin rgb_reg = 3'b111; end
            18'b101011001011010001: begin rgb_reg = 3'b111; end
            18'b101011001011010010: begin rgb_reg = 3'b111; end
            18'b101011001011010011: begin rgb_reg = 3'b111; end
            18'b101011001011010100: begin rgb_reg = 3'b111; end
            18'b101011001011011001: begin rgb_reg = 3'b111; end
            18'b101011001011011010: begin rgb_reg = 3'b111; end
            18'b101011001011100001: begin rgb_reg = 3'b111; end
            18'b101011001011100010: begin rgb_reg = 3'b111; end
            18'b101011001011100101: begin rgb_reg = 3'b111; end
            18'b101011001011100110: begin rgb_reg = 3'b111; end
            18'b101011001011100111: begin rgb_reg = 3'b111; end
            18'b101011001011101000: begin rgb_reg = 3'b111; end
            18'b101011001011101011: begin rgb_reg = 3'b111; end
            18'b101011001011101100: begin rgb_reg = 3'b111; end
            18'b101011001011111101: begin rgb_reg = 3'b111; end
            18'b101011001011111110: begin rgb_reg = 3'b111; end
            18'b101011001100000001: begin rgb_reg = 3'b111; end
            18'b101011001100000010: begin rgb_reg = 3'b111; end
            18'b101011001100000101: begin rgb_reg = 3'b111; end
            18'b101011001100000110: begin rgb_reg = 3'b111; end
            18'b101011001100001001: begin rgb_reg = 3'b111; end
            18'b101011001100001010: begin rgb_reg = 3'b111; end
            18'b101011001100001101: begin rgb_reg = 3'b111; end
            18'b101011001100001110: begin rgb_reg = 3'b111; end
            18'b101011001100010101: begin rgb_reg = 3'b111; end
            18'b101011001100010110: begin rgb_reg = 3'b111; end
            18'b101011001100011011: begin rgb_reg = 3'b111; end
            18'b101011001100011100: begin rgb_reg = 3'b111; end
            18'b101011001100011101: begin rgb_reg = 3'b111; end
            18'b101011001100011110: begin rgb_reg = 3'b111; end
            18'b101011001100011111: begin rgb_reg = 3'b111; end
            18'b101011001100100000: begin rgb_reg = 3'b111; end
            18'b101011001100100101: begin rgb_reg = 3'b111; end
            18'b101011001100100110: begin rgb_reg = 3'b111; end
            18'b101011001100100111: begin rgb_reg = 3'b111; end
            18'b101011001100101000: begin rgb_reg = 3'b111; end
            18'b101011001100101011: begin rgb_reg = 3'b111; end
            18'b101011001100101100: begin rgb_reg = 3'b111; end
            18'b101011001100110011: begin rgb_reg = 3'b111; end
            18'b101011001100110100: begin rgb_reg = 3'b111; end
            18'b101011001100110101: begin rgb_reg = 3'b111; end
            18'b101011001100110110: begin rgb_reg = 3'b111; end
            18'b101011001100110111: begin rgb_reg = 3'b111; end
            18'b101011001100111000: begin rgb_reg = 3'b111; end
            18'b101011001100111001: begin rgb_reg = 3'b111; end
            18'b101011001100111010: begin rgb_reg = 3'b111; end
            18'b101011001100111111: begin rgb_reg = 3'b111; end
            18'b101011001101000000: begin rgb_reg = 3'b111; end
            18'b101011001101000001: begin rgb_reg = 3'b111; end
            18'b101011001101000010: begin rgb_reg = 3'b111; end
            18'b101011001101000011: begin rgb_reg = 3'b111; end
            18'b101011001101000100: begin rgb_reg = 3'b111; end
            18'b101011001101001011: begin rgb_reg = 3'b111; end
            18'b101011001101001100: begin rgb_reg = 3'b111; end
            18'b101011001101010001: begin rgb_reg = 3'b111; end
            18'b101011001101010010: begin rgb_reg = 3'b111; end
            18'b101011001101010101: begin rgb_reg = 3'b111; end
            18'b101011001101010110: begin rgb_reg = 3'b111; end
            18'b101011001101010111: begin rgb_reg = 3'b111; end
            18'b101011001101011000: begin rgb_reg = 3'b111; end
            18'b101011001101011101: begin rgb_reg = 3'b111; end
            18'b101011001101011110: begin rgb_reg = 3'b111; end
            18'b101011001101100011: begin rgb_reg = 3'b111; end
            18'b101011001101100100: begin rgb_reg = 3'b111; end
            18'b101011001101100101: begin rgb_reg = 3'b111; end
            18'b101011001101100110: begin rgb_reg = 3'b111; end
            18'b101011001101100111: begin rgb_reg = 3'b111; end
            18'b101011001101101000: begin rgb_reg = 3'b111; end
            18'b101011001101101101: begin rgb_reg = 3'b111; end
            18'b101011001101101110: begin rgb_reg = 3'b111; end
            18'b101011001101101111: begin rgb_reg = 3'b111; end
            18'b101011001101110000: begin rgb_reg = 3'b111; end
            18'b101011001101110001: begin rgb_reg = 3'b111; end
            18'b101011001101110010: begin rgb_reg = 3'b111; end
            18'b101011001101110011: begin rgb_reg = 3'b111; end
            18'b101011001101110100: begin rgb_reg = 3'b111; end
            18'b101011010010001001: begin rgb_reg = 3'b111; end
            18'b101011010010001010: begin rgb_reg = 3'b111; end
            18'b101011010010001101: begin rgb_reg = 3'b111; end
            18'b101011010010001110: begin rgb_reg = 3'b111; end
            18'b101011010010010001: begin rgb_reg = 3'b111; end
            18'b101011010010010010: begin rgb_reg = 3'b111; end
            18'b101011010010010111: begin rgb_reg = 3'b111; end
            18'b101011010010011000: begin rgb_reg = 3'b111; end
            18'b101011010010011001: begin rgb_reg = 3'b111; end
            18'b101011010010011010: begin rgb_reg = 3'b111; end
            18'b101011010010011011: begin rgb_reg = 3'b111; end
            18'b101011010010011100: begin rgb_reg = 3'b111; end
            18'b101011010010100011: begin rgb_reg = 3'b111; end
            18'b101011010010100100: begin rgb_reg = 3'b111; end
            18'b101011010010101001: begin rgb_reg = 3'b111; end
            18'b101011010010101010: begin rgb_reg = 3'b111; end
            18'b101011010010101101: begin rgb_reg = 3'b111; end
            18'b101011010010101110: begin rgb_reg = 3'b111; end
            18'b101011010010101111: begin rgb_reg = 3'b111; end
            18'b101011010010110000: begin rgb_reg = 3'b111; end
            18'b101011010010110111: begin rgb_reg = 3'b111; end
            18'b101011010010111000: begin rgb_reg = 3'b111; end
            18'b101011010010111001: begin rgb_reg = 3'b111; end
            18'b101011010010111010: begin rgb_reg = 3'b111; end
            18'b101011010010111011: begin rgb_reg = 3'b111; end
            18'b101011010010111100: begin rgb_reg = 3'b111; end
            18'b101011010011000001: begin rgb_reg = 3'b111; end
            18'b101011010011000010: begin rgb_reg = 3'b111; end
            18'b101011010011000101: begin rgb_reg = 3'b111; end
            18'b101011010011000110: begin rgb_reg = 3'b111; end
            18'b101011010011000111: begin rgb_reg = 3'b111; end
            18'b101011010011001000: begin rgb_reg = 3'b111; end
            18'b101011010011001101: begin rgb_reg = 3'b111; end
            18'b101011010011001110: begin rgb_reg = 3'b111; end
            18'b101011010011010001: begin rgb_reg = 3'b111; end
            18'b101011010011010010: begin rgb_reg = 3'b111; end
            18'b101011010011010011: begin rgb_reg = 3'b111; end
            18'b101011010011010100: begin rgb_reg = 3'b111; end
            18'b101011010011011001: begin rgb_reg = 3'b111; end
            18'b101011010011011010: begin rgb_reg = 3'b111; end
            18'b101011010011100001: begin rgb_reg = 3'b111; end
            18'b101011010011100010: begin rgb_reg = 3'b111; end
            18'b101011010011100101: begin rgb_reg = 3'b111; end
            18'b101011010011100110: begin rgb_reg = 3'b111; end
            18'b101011010011100111: begin rgb_reg = 3'b111; end
            18'b101011010011101000: begin rgb_reg = 3'b111; end
            18'b101011010011101011: begin rgb_reg = 3'b111; end
            18'b101011010011101100: begin rgb_reg = 3'b111; end
            18'b101011010011111101: begin rgb_reg = 3'b111; end
            18'b101011010011111110: begin rgb_reg = 3'b111; end
            18'b101011010100000001: begin rgb_reg = 3'b111; end
            18'b101011010100000010: begin rgb_reg = 3'b111; end
            18'b101011010100000101: begin rgb_reg = 3'b111; end
            18'b101011010100000110: begin rgb_reg = 3'b111; end
            18'b101011010100001001: begin rgb_reg = 3'b111; end
            18'b101011010100001010: begin rgb_reg = 3'b111; end
            18'b101011010100001101: begin rgb_reg = 3'b111; end
            18'b101011010100001110: begin rgb_reg = 3'b111; end
            18'b101011010100010101: begin rgb_reg = 3'b111; end
            18'b101011010100010110: begin rgb_reg = 3'b111; end
            18'b101011010100011011: begin rgb_reg = 3'b111; end
            18'b101011010100011100: begin rgb_reg = 3'b111; end
            18'b101011010100011101: begin rgb_reg = 3'b111; end
            18'b101011010100011110: begin rgb_reg = 3'b111; end
            18'b101011010100011111: begin rgb_reg = 3'b111; end
            18'b101011010100100000: begin rgb_reg = 3'b111; end
            18'b101011010100100101: begin rgb_reg = 3'b111; end
            18'b101011010100100110: begin rgb_reg = 3'b111; end
            18'b101011010100100111: begin rgb_reg = 3'b111; end
            18'b101011010100101000: begin rgb_reg = 3'b111; end
            18'b101011010100101011: begin rgb_reg = 3'b111; end
            18'b101011010100101100: begin rgb_reg = 3'b111; end
            18'b101011010100110011: begin rgb_reg = 3'b111; end
            18'b101011010100110100: begin rgb_reg = 3'b111; end
            18'b101011010100110101: begin rgb_reg = 3'b111; end
            18'b101011010100110110: begin rgb_reg = 3'b111; end
            18'b101011010100110111: begin rgb_reg = 3'b111; end
            18'b101011010100111000: begin rgb_reg = 3'b111; end
            18'b101011010100111001: begin rgb_reg = 3'b111; end
            18'b101011010100111010: begin rgb_reg = 3'b111; end
            18'b101011010100111111: begin rgb_reg = 3'b111; end
            18'b101011010101000000: begin rgb_reg = 3'b111; end
            18'b101011010101000001: begin rgb_reg = 3'b111; end
            18'b101011010101000010: begin rgb_reg = 3'b111; end
            18'b101011010101000011: begin rgb_reg = 3'b111; end
            18'b101011010101000100: begin rgb_reg = 3'b111; end
            18'b101011010101001011: begin rgb_reg = 3'b111; end
            18'b101011010101001100: begin rgb_reg = 3'b111; end
            18'b101011010101010001: begin rgb_reg = 3'b111; end
            18'b101011010101010010: begin rgb_reg = 3'b111; end
            18'b101011010101010101: begin rgb_reg = 3'b111; end
            18'b101011010101010110: begin rgb_reg = 3'b111; end
            18'b101011010101010111: begin rgb_reg = 3'b111; end
            18'b101011010101011000: begin rgb_reg = 3'b111; end
            18'b101011010101011101: begin rgb_reg = 3'b111; end
            18'b101011010101011110: begin rgb_reg = 3'b111; end
            18'b101011010101100011: begin rgb_reg = 3'b111; end
            18'b101011010101100100: begin rgb_reg = 3'b111; end
            18'b101011010101100101: begin rgb_reg = 3'b111; end
            18'b101011010101100110: begin rgb_reg = 3'b111; end
            18'b101011010101100111: begin rgb_reg = 3'b111; end
            18'b101011010101101000: begin rgb_reg = 3'b111; end
            18'b101011010101101101: begin rgb_reg = 3'b111; end
            18'b101011010101101110: begin rgb_reg = 3'b111; end
            18'b101011010101101111: begin rgb_reg = 3'b111; end
            18'b101011010101110000: begin rgb_reg = 3'b111; end
            18'b101011010101110001: begin rgb_reg = 3'b111; end
            18'b101011010101110010: begin rgb_reg = 3'b111; end
            18'b101011010101110011: begin rgb_reg = 3'b111; end
            18'b101011010101110100: begin rgb_reg = 3'b111; end
            18'b101011011010001001: begin rgb_reg = 3'b111; end
            18'b101011011010001010: begin rgb_reg = 3'b111; end
            18'b101011011010001111: begin rgb_reg = 3'b111; end
            18'b101011011010010000: begin rgb_reg = 3'b111; end
            18'b101011011010010001: begin rgb_reg = 3'b111; end
            18'b101011011010010010: begin rgb_reg = 3'b111; end
            18'b101011011010011101: begin rgb_reg = 3'b111; end
            18'b101011011010011110: begin rgb_reg = 3'b111; end
            18'b101011011010100011: begin rgb_reg = 3'b111; end
            18'b101011011010100100: begin rgb_reg = 3'b111; end
            18'b101011011010101001: begin rgb_reg = 3'b111; end
            18'b101011011010101010: begin rgb_reg = 3'b111; end
            18'b101011011010101011: begin rgb_reg = 3'b111; end
            18'b101011011010101100: begin rgb_reg = 3'b111; end
            18'b101011011010110001: begin rgb_reg = 3'b111; end
            18'b101011011010110010: begin rgb_reg = 3'b111; end
            18'b101011011010111101: begin rgb_reg = 3'b111; end
            18'b101011011010111110: begin rgb_reg = 3'b111; end
            18'b101011011011000001: begin rgb_reg = 3'b111; end
            18'b101011011011000010: begin rgb_reg = 3'b111; end
            18'b101011011011000011: begin rgb_reg = 3'b111; end
            18'b101011011011000100: begin rgb_reg = 3'b111; end
            18'b101011011011001001: begin rgb_reg = 3'b111; end
            18'b101011011011001010: begin rgb_reg = 3'b111; end
            18'b101011011011001101: begin rgb_reg = 3'b111; end
            18'b101011011011001110: begin rgb_reg = 3'b111; end
            18'b101011011011001111: begin rgb_reg = 3'b111; end
            18'b101011011011010000: begin rgb_reg = 3'b111; end
            18'b101011011011010101: begin rgb_reg = 3'b111; end
            18'b101011011011010110: begin rgb_reg = 3'b111; end
            18'b101011011011011001: begin rgb_reg = 3'b111; end
            18'b101011011011011010: begin rgb_reg = 3'b111; end
            18'b101011011011100001: begin rgb_reg = 3'b111; end
            18'b101011011011100010: begin rgb_reg = 3'b111; end
            18'b101011011011100101: begin rgb_reg = 3'b111; end
            18'b101011011011100110: begin rgb_reg = 3'b111; end
            18'b101011011011101001: begin rgb_reg = 3'b111; end
            18'b101011011011101010: begin rgb_reg = 3'b111; end
            18'b101011011011101101: begin rgb_reg = 3'b111; end
            18'b101011011011101110: begin rgb_reg = 3'b111; end
            18'b101011011011111101: begin rgb_reg = 3'b111; end
            18'b101011011011111110: begin rgb_reg = 3'b111; end
            18'b101011011100000011: begin rgb_reg = 3'b111; end
            18'b101011011100000100: begin rgb_reg = 3'b111; end
            18'b101011011100000101: begin rgb_reg = 3'b111; end
            18'b101011011100000110: begin rgb_reg = 3'b111; end
            18'b101011011100001001: begin rgb_reg = 3'b111; end
            18'b101011011100001010: begin rgb_reg = 3'b111; end
            18'b101011011100001101: begin rgb_reg = 3'b111; end
            18'b101011011100001110: begin rgb_reg = 3'b111; end
            18'b101011011100010101: begin rgb_reg = 3'b111; end
            18'b101011011100010110: begin rgb_reg = 3'b111; end
            18'b101011011100011001: begin rgb_reg = 3'b111; end
            18'b101011011100011010: begin rgb_reg = 3'b111; end
            18'b101011011100100001: begin rgb_reg = 3'b111; end
            18'b101011011100100010: begin rgb_reg = 3'b111; end
            18'b101011011100100101: begin rgb_reg = 3'b111; end
            18'b101011011100100110: begin rgb_reg = 3'b111; end
            18'b101011011100101001: begin rgb_reg = 3'b111; end
            18'b101011011100101010: begin rgb_reg = 3'b111; end
            18'b101011011100101101: begin rgb_reg = 3'b111; end
            18'b101011011100101110: begin rgb_reg = 3'b111; end
            18'b101011011100110001: begin rgb_reg = 3'b111; end
            18'b101011011100110010: begin rgb_reg = 3'b111; end
            18'b101011011101000101: begin rgb_reg = 3'b111; end
            18'b101011011101000110: begin rgb_reg = 3'b111; end
            18'b101011011101001011: begin rgb_reg = 3'b111; end
            18'b101011011101001100: begin rgb_reg = 3'b111; end
            18'b101011011101010001: begin rgb_reg = 3'b111; end
            18'b101011011101010010: begin rgb_reg = 3'b111; end
            18'b101011011101010011: begin rgb_reg = 3'b111; end
            18'b101011011101010100: begin rgb_reg = 3'b111; end
            18'b101011011101011001: begin rgb_reg = 3'b111; end
            18'b101011011101011010: begin rgb_reg = 3'b111; end
            18'b101011011101011101: begin rgb_reg = 3'b111; end
            18'b101011011101011110: begin rgb_reg = 3'b111; end
            18'b101011011101100001: begin rgb_reg = 3'b111; end
            18'b101011011101100010: begin rgb_reg = 3'b111; end
            18'b101011011101101001: begin rgb_reg = 3'b111; end
            18'b101011011101101010: begin rgb_reg = 3'b111; end
            18'b101011011101101101: begin rgb_reg = 3'b111; end
            18'b101011011101101110: begin rgb_reg = 3'b111; end
            18'b101011011101110101: begin rgb_reg = 3'b111; end
            18'b101011011101110110: begin rgb_reg = 3'b111; end
            18'b101011100010001001: begin rgb_reg = 3'b111; end
            18'b101011100010001010: begin rgb_reg = 3'b111; end
            18'b101011100010001111: begin rgb_reg = 3'b111; end
            18'b101011100010010000: begin rgb_reg = 3'b111; end
            18'b101011100010010001: begin rgb_reg = 3'b111; end
            18'b101011100010010010: begin rgb_reg = 3'b111; end
            18'b101011100010011101: begin rgb_reg = 3'b111; end
            18'b101011100010011110: begin rgb_reg = 3'b111; end
            18'b101011100010100011: begin rgb_reg = 3'b111; end
            18'b101011100010100100: begin rgb_reg = 3'b111; end
            18'b101011100010101001: begin rgb_reg = 3'b111; end
            18'b101011100010101010: begin rgb_reg = 3'b111; end
            18'b101011100010101011: begin rgb_reg = 3'b111; end
            18'b101011100010101100: begin rgb_reg = 3'b111; end
            18'b101011100010110001: begin rgb_reg = 3'b111; end
            18'b101011100010110010: begin rgb_reg = 3'b111; end
            18'b101011100010111101: begin rgb_reg = 3'b111; end
            18'b101011100010111110: begin rgb_reg = 3'b111; end
            18'b101011100011000001: begin rgb_reg = 3'b111; end
            18'b101011100011000010: begin rgb_reg = 3'b111; end
            18'b101011100011000011: begin rgb_reg = 3'b111; end
            18'b101011100011000100: begin rgb_reg = 3'b111; end
            18'b101011100011001001: begin rgb_reg = 3'b111; end
            18'b101011100011001010: begin rgb_reg = 3'b111; end
            18'b101011100011001101: begin rgb_reg = 3'b111; end
            18'b101011100011001110: begin rgb_reg = 3'b111; end
            18'b101011100011001111: begin rgb_reg = 3'b111; end
            18'b101011100011010000: begin rgb_reg = 3'b111; end
            18'b101011100011010101: begin rgb_reg = 3'b111; end
            18'b101011100011010110: begin rgb_reg = 3'b111; end
            18'b101011100011011001: begin rgb_reg = 3'b111; end
            18'b101011100011011010: begin rgb_reg = 3'b111; end
            18'b101011100011100001: begin rgb_reg = 3'b111; end
            18'b101011100011100010: begin rgb_reg = 3'b111; end
            18'b101011100011100101: begin rgb_reg = 3'b111; end
            18'b101011100011100110: begin rgb_reg = 3'b111; end
            18'b101011100011101001: begin rgb_reg = 3'b111; end
            18'b101011100011101010: begin rgb_reg = 3'b111; end
            18'b101011100011101101: begin rgb_reg = 3'b111; end
            18'b101011100011101110: begin rgb_reg = 3'b111; end
            18'b101011100011111101: begin rgb_reg = 3'b111; end
            18'b101011100011111110: begin rgb_reg = 3'b111; end
            18'b101011100100000011: begin rgb_reg = 3'b111; end
            18'b101011100100000100: begin rgb_reg = 3'b111; end
            18'b101011100100000101: begin rgb_reg = 3'b111; end
            18'b101011100100000110: begin rgb_reg = 3'b111; end
            18'b101011100100001001: begin rgb_reg = 3'b111; end
            18'b101011100100001010: begin rgb_reg = 3'b111; end
            18'b101011100100001101: begin rgb_reg = 3'b111; end
            18'b101011100100001110: begin rgb_reg = 3'b111; end
            18'b101011100100010101: begin rgb_reg = 3'b111; end
            18'b101011100100010110: begin rgb_reg = 3'b111; end
            18'b101011100100011001: begin rgb_reg = 3'b111; end
            18'b101011100100011010: begin rgb_reg = 3'b111; end
            18'b101011100100100001: begin rgb_reg = 3'b111; end
            18'b101011100100100010: begin rgb_reg = 3'b111; end
            18'b101011100100100101: begin rgb_reg = 3'b111; end
            18'b101011100100100110: begin rgb_reg = 3'b111; end
            18'b101011100100101001: begin rgb_reg = 3'b111; end
            18'b101011100100101010: begin rgb_reg = 3'b111; end
            18'b101011100100101101: begin rgb_reg = 3'b111; end
            18'b101011100100101110: begin rgb_reg = 3'b111; end
            18'b101011100100110001: begin rgb_reg = 3'b111; end
            18'b101011100100110010: begin rgb_reg = 3'b111; end
            18'b101011100101000101: begin rgb_reg = 3'b111; end
            18'b101011100101000110: begin rgb_reg = 3'b111; end
            18'b101011100101001011: begin rgb_reg = 3'b111; end
            18'b101011100101001100: begin rgb_reg = 3'b111; end
            18'b101011100101010001: begin rgb_reg = 3'b111; end
            18'b101011100101010010: begin rgb_reg = 3'b111; end
            18'b101011100101010011: begin rgb_reg = 3'b111; end
            18'b101011100101010100: begin rgb_reg = 3'b111; end
            18'b101011100101011001: begin rgb_reg = 3'b111; end
            18'b101011100101011010: begin rgb_reg = 3'b111; end
            18'b101011100101011101: begin rgb_reg = 3'b111; end
            18'b101011100101011110: begin rgb_reg = 3'b111; end
            18'b101011100101100001: begin rgb_reg = 3'b111; end
            18'b101011100101100010: begin rgb_reg = 3'b111; end
            18'b101011100101101001: begin rgb_reg = 3'b111; end
            18'b101011100101101010: begin rgb_reg = 3'b111; end
            18'b101011100101101101: begin rgb_reg = 3'b111; end
            18'b101011100101101110: begin rgb_reg = 3'b111; end
            18'b101011100101110101: begin rgb_reg = 3'b111; end
            18'b101011100101110110: begin rgb_reg = 3'b111; end
            18'b101011101010001001: begin rgb_reg = 3'b111; end
            18'b101011101010001010: begin rgb_reg = 3'b111; end
            18'b101011101010010001: begin rgb_reg = 3'b111; end
            18'b101011101010010010: begin rgb_reg = 3'b111; end
            18'b101011101010010111: begin rgb_reg = 3'b111; end
            18'b101011101010011000: begin rgb_reg = 3'b111; end
            18'b101011101010011001: begin rgb_reg = 3'b111; end
            18'b101011101010011010: begin rgb_reg = 3'b111; end
            18'b101011101010011011: begin rgb_reg = 3'b111; end
            18'b101011101010011100: begin rgb_reg = 3'b111; end
            18'b101011101010011101: begin rgb_reg = 3'b111; end
            18'b101011101010011110: begin rgb_reg = 3'b111; end
            18'b101011101010100011: begin rgb_reg = 3'b111; end
            18'b101011101010100100: begin rgb_reg = 3'b111; end
            18'b101011101010101001: begin rgb_reg = 3'b111; end
            18'b101011101010101010: begin rgb_reg = 3'b111; end
            18'b101011101010110001: begin rgb_reg = 3'b111; end
            18'b101011101010110010: begin rgb_reg = 3'b111; end
            18'b101011101010110111: begin rgb_reg = 3'b111; end
            18'b101011101010111000: begin rgb_reg = 3'b111; end
            18'b101011101010111001: begin rgb_reg = 3'b111; end
            18'b101011101010111010: begin rgb_reg = 3'b111; end
            18'b101011101010111011: begin rgb_reg = 3'b111; end
            18'b101011101010111100: begin rgb_reg = 3'b111; end
            18'b101011101010111101: begin rgb_reg = 3'b111; end
            18'b101011101010111110: begin rgb_reg = 3'b111; end
            18'b101011101011000001: begin rgb_reg = 3'b111; end
            18'b101011101011000010: begin rgb_reg = 3'b111; end
            18'b101011101011001001: begin rgb_reg = 3'b111; end
            18'b101011101011001010: begin rgb_reg = 3'b111; end
            18'b101011101011001101: begin rgb_reg = 3'b111; end
            18'b101011101011001110: begin rgb_reg = 3'b111; end
            18'b101011101011010101: begin rgb_reg = 3'b111; end
            18'b101011101011010110: begin rgb_reg = 3'b111; end
            18'b101011101011011001: begin rgb_reg = 3'b111; end
            18'b101011101011011010: begin rgb_reg = 3'b111; end
            18'b101011101011100001: begin rgb_reg = 3'b111; end
            18'b101011101011100010: begin rgb_reg = 3'b111; end
            18'b101011101011100101: begin rgb_reg = 3'b111; end
            18'b101011101011100110: begin rgb_reg = 3'b111; end
            18'b101011101011101001: begin rgb_reg = 3'b111; end
            18'b101011101011101010: begin rgb_reg = 3'b111; end
            18'b101011101011101101: begin rgb_reg = 3'b111; end
            18'b101011101011101110: begin rgb_reg = 3'b111; end
            18'b101011101011111101: begin rgb_reg = 3'b111; end
            18'b101011101011111110: begin rgb_reg = 3'b111; end
            18'b101011101100000101: begin rgb_reg = 3'b111; end
            18'b101011101100000110: begin rgb_reg = 3'b111; end
            18'b101011101100001001: begin rgb_reg = 3'b111; end
            18'b101011101100001010: begin rgb_reg = 3'b111; end
            18'b101011101100001101: begin rgb_reg = 3'b111; end
            18'b101011101100001110: begin rgb_reg = 3'b111; end
            18'b101011101100010101: begin rgb_reg = 3'b111; end
            18'b101011101100010110: begin rgb_reg = 3'b111; end
            18'b101011101100011001: begin rgb_reg = 3'b111; end
            18'b101011101100011010: begin rgb_reg = 3'b111; end
            18'b101011101100100001: begin rgb_reg = 3'b111; end
            18'b101011101100100010: begin rgb_reg = 3'b111; end
            18'b101011101100100101: begin rgb_reg = 3'b111; end
            18'b101011101100100110: begin rgb_reg = 3'b111; end
            18'b101011101100101001: begin rgb_reg = 3'b111; end
            18'b101011101100101010: begin rgb_reg = 3'b111; end
            18'b101011101100101101: begin rgb_reg = 3'b111; end
            18'b101011101100101110: begin rgb_reg = 3'b111; end
            18'b101011101100110011: begin rgb_reg = 3'b111; end
            18'b101011101100110100: begin rgb_reg = 3'b111; end
            18'b101011101100110101: begin rgb_reg = 3'b111; end
            18'b101011101100110110: begin rgb_reg = 3'b111; end
            18'b101011101100110111: begin rgb_reg = 3'b111; end
            18'b101011101100111000: begin rgb_reg = 3'b111; end
            18'b101011101100111111: begin rgb_reg = 3'b111; end
            18'b101011101101000000: begin rgb_reg = 3'b111; end
            18'b101011101101000001: begin rgb_reg = 3'b111; end
            18'b101011101101000010: begin rgb_reg = 3'b111; end
            18'b101011101101000011: begin rgb_reg = 3'b111; end
            18'b101011101101000100: begin rgb_reg = 3'b111; end
            18'b101011101101000101: begin rgb_reg = 3'b111; end
            18'b101011101101000110: begin rgb_reg = 3'b111; end
            18'b101011101101001011: begin rgb_reg = 3'b111; end
            18'b101011101101001100: begin rgb_reg = 3'b111; end
            18'b101011101101010001: begin rgb_reg = 3'b111; end
            18'b101011101101010010: begin rgb_reg = 3'b111; end
            18'b101011101101011001: begin rgb_reg = 3'b111; end
            18'b101011101101011010: begin rgb_reg = 3'b111; end
            18'b101011101101011101: begin rgb_reg = 3'b111; end
            18'b101011101101011110: begin rgb_reg = 3'b111; end
            18'b101011101101100001: begin rgb_reg = 3'b111; end
            18'b101011101101100010: begin rgb_reg = 3'b111; end
            18'b101011101101100011: begin rgb_reg = 3'b111; end
            18'b101011101101100100: begin rgb_reg = 3'b111; end
            18'b101011101101100101: begin rgb_reg = 3'b111; end
            18'b101011101101100110: begin rgb_reg = 3'b111; end
            18'b101011101101100111: begin rgb_reg = 3'b111; end
            18'b101011101101101000: begin rgb_reg = 3'b111; end
            18'b101011101101101001: begin rgb_reg = 3'b111; end
            18'b101011101101101010: begin rgb_reg = 3'b111; end
            18'b101011101101101101: begin rgb_reg = 3'b111; end
            18'b101011101101101110: begin rgb_reg = 3'b111; end
            18'b101011101101110101: begin rgb_reg = 3'b111; end
            18'b101011101101110110: begin rgb_reg = 3'b111; end
            18'b101011110010001001: begin rgb_reg = 3'b111; end
            18'b101011110010001010: begin rgb_reg = 3'b111; end
            18'b101011110010010001: begin rgb_reg = 3'b111; end
            18'b101011110010010010: begin rgb_reg = 3'b111; end
            18'b101011110010010111: begin rgb_reg = 3'b111; end
            18'b101011110010011000: begin rgb_reg = 3'b111; end
            18'b101011110010011001: begin rgb_reg = 3'b111; end
            18'b101011110010011010: begin rgb_reg = 3'b111; end
            18'b101011110010011011: begin rgb_reg = 3'b111; end
            18'b101011110010011100: begin rgb_reg = 3'b111; end
            18'b101011110010011101: begin rgb_reg = 3'b111; end
            18'b101011110010011110: begin rgb_reg = 3'b111; end
            18'b101011110010100011: begin rgb_reg = 3'b111; end
            18'b101011110010100100: begin rgb_reg = 3'b111; end
            18'b101011110010101001: begin rgb_reg = 3'b111; end
            18'b101011110010101010: begin rgb_reg = 3'b111; end
            18'b101011110010110001: begin rgb_reg = 3'b111; end
            18'b101011110010110010: begin rgb_reg = 3'b111; end
            18'b101011110010110111: begin rgb_reg = 3'b111; end
            18'b101011110010111000: begin rgb_reg = 3'b111; end
            18'b101011110010111001: begin rgb_reg = 3'b111; end
            18'b101011110010111010: begin rgb_reg = 3'b111; end
            18'b101011110010111011: begin rgb_reg = 3'b111; end
            18'b101011110010111100: begin rgb_reg = 3'b111; end
            18'b101011110010111101: begin rgb_reg = 3'b111; end
            18'b101011110010111110: begin rgb_reg = 3'b111; end
            18'b101011110011000001: begin rgb_reg = 3'b111; end
            18'b101011110011000010: begin rgb_reg = 3'b111; end
            18'b101011110011001001: begin rgb_reg = 3'b111; end
            18'b101011110011001010: begin rgb_reg = 3'b111; end
            18'b101011110011001101: begin rgb_reg = 3'b111; end
            18'b101011110011001110: begin rgb_reg = 3'b111; end
            18'b101011110011010101: begin rgb_reg = 3'b111; end
            18'b101011110011010110: begin rgb_reg = 3'b111; end
            18'b101011110011011001: begin rgb_reg = 3'b111; end
            18'b101011110011011010: begin rgb_reg = 3'b111; end
            18'b101011110011100001: begin rgb_reg = 3'b111; end
            18'b101011110011100010: begin rgb_reg = 3'b111; end
            18'b101011110011100101: begin rgb_reg = 3'b111; end
            18'b101011110011100110: begin rgb_reg = 3'b111; end
            18'b101011110011101001: begin rgb_reg = 3'b111; end
            18'b101011110011101010: begin rgb_reg = 3'b111; end
            18'b101011110011101101: begin rgb_reg = 3'b111; end
            18'b101011110011101110: begin rgb_reg = 3'b111; end
            18'b101011110011111101: begin rgb_reg = 3'b111; end
            18'b101011110011111110: begin rgb_reg = 3'b111; end
            18'b101011110100000101: begin rgb_reg = 3'b111; end
            18'b101011110100000110: begin rgb_reg = 3'b111; end
            18'b101011110100001001: begin rgb_reg = 3'b111; end
            18'b101011110100001010: begin rgb_reg = 3'b111; end
            18'b101011110100001101: begin rgb_reg = 3'b111; end
            18'b101011110100001110: begin rgb_reg = 3'b111; end
            18'b101011110100010101: begin rgb_reg = 3'b111; end
            18'b101011110100010110: begin rgb_reg = 3'b111; end
            18'b101011110100011001: begin rgb_reg = 3'b111; end
            18'b101011110100011010: begin rgb_reg = 3'b111; end
            18'b101011110100100001: begin rgb_reg = 3'b111; end
            18'b101011110100100010: begin rgb_reg = 3'b111; end
            18'b101011110100100101: begin rgb_reg = 3'b111; end
            18'b101011110100100110: begin rgb_reg = 3'b111; end
            18'b101011110100101001: begin rgb_reg = 3'b111; end
            18'b101011110100101010: begin rgb_reg = 3'b111; end
            18'b101011110100101101: begin rgb_reg = 3'b111; end
            18'b101011110100101110: begin rgb_reg = 3'b111; end
            18'b101011110100110011: begin rgb_reg = 3'b111; end
            18'b101011110100110100: begin rgb_reg = 3'b111; end
            18'b101011110100110101: begin rgb_reg = 3'b111; end
            18'b101011110100110110: begin rgb_reg = 3'b111; end
            18'b101011110100110111: begin rgb_reg = 3'b111; end
            18'b101011110100111000: begin rgb_reg = 3'b111; end
            18'b101011110100111111: begin rgb_reg = 3'b111; end
            18'b101011110101000000: begin rgb_reg = 3'b111; end
            18'b101011110101000001: begin rgb_reg = 3'b111; end
            18'b101011110101000010: begin rgb_reg = 3'b111; end
            18'b101011110101000011: begin rgb_reg = 3'b111; end
            18'b101011110101000100: begin rgb_reg = 3'b111; end
            18'b101011110101000101: begin rgb_reg = 3'b111; end
            18'b101011110101000110: begin rgb_reg = 3'b111; end
            18'b101011110101001011: begin rgb_reg = 3'b111; end
            18'b101011110101001100: begin rgb_reg = 3'b111; end
            18'b101011110101010001: begin rgb_reg = 3'b111; end
            18'b101011110101010010: begin rgb_reg = 3'b111; end
            18'b101011110101011001: begin rgb_reg = 3'b111; end
            18'b101011110101011010: begin rgb_reg = 3'b111; end
            18'b101011110101011101: begin rgb_reg = 3'b111; end
            18'b101011110101011110: begin rgb_reg = 3'b111; end
            18'b101011110101100001: begin rgb_reg = 3'b111; end
            18'b101011110101100010: begin rgb_reg = 3'b111; end
            18'b101011110101100011: begin rgb_reg = 3'b111; end
            18'b101011110101100100: begin rgb_reg = 3'b111; end
            18'b101011110101100101: begin rgb_reg = 3'b111; end
            18'b101011110101100110: begin rgb_reg = 3'b111; end
            18'b101011110101100111: begin rgb_reg = 3'b111; end
            18'b101011110101101000: begin rgb_reg = 3'b111; end
            18'b101011110101101001: begin rgb_reg = 3'b111; end
            18'b101011110101101010: begin rgb_reg = 3'b111; end
            18'b101011110101101101: begin rgb_reg = 3'b111; end
            18'b101011110101101110: begin rgb_reg = 3'b111; end
            18'b101011110101110101: begin rgb_reg = 3'b111; end
            18'b101011110101110110: begin rgb_reg = 3'b111; end
            18'b101011111010001001: begin rgb_reg = 3'b111; end
            18'b101011111010001010: begin rgb_reg = 3'b111; end
            18'b101011111010010001: begin rgb_reg = 3'b111; end
            18'b101011111010010010: begin rgb_reg = 3'b111; end
            18'b101011111010010101: begin rgb_reg = 3'b111; end
            18'b101011111010010110: begin rgb_reg = 3'b111; end
            18'b101011111010011101: begin rgb_reg = 3'b111; end
            18'b101011111010011110: begin rgb_reg = 3'b111; end
            18'b101011111010100011: begin rgb_reg = 3'b111; end
            18'b101011111010100100: begin rgb_reg = 3'b111; end
            18'b101011111010101001: begin rgb_reg = 3'b111; end
            18'b101011111010101010: begin rgb_reg = 3'b111; end
            18'b101011111010110001: begin rgb_reg = 3'b111; end
            18'b101011111010110010: begin rgb_reg = 3'b111; end
            18'b101011111010110101: begin rgb_reg = 3'b111; end
            18'b101011111010110110: begin rgb_reg = 3'b111; end
            18'b101011111010111101: begin rgb_reg = 3'b111; end
            18'b101011111010111110: begin rgb_reg = 3'b111; end
            18'b101011111011000001: begin rgb_reg = 3'b111; end
            18'b101011111011000010: begin rgb_reg = 3'b111; end
            18'b101011111011000011: begin rgb_reg = 3'b111; end
            18'b101011111011000100: begin rgb_reg = 3'b111; end
            18'b101011111011000101: begin rgb_reg = 3'b111; end
            18'b101011111011000110: begin rgb_reg = 3'b111; end
            18'b101011111011000111: begin rgb_reg = 3'b111; end
            18'b101011111011001000: begin rgb_reg = 3'b111; end
            18'b101011111011001101: begin rgb_reg = 3'b111; end
            18'b101011111011001110: begin rgb_reg = 3'b111; end
            18'b101011111011010101: begin rgb_reg = 3'b111; end
            18'b101011111011010110: begin rgb_reg = 3'b111; end
            18'b101011111011011001: begin rgb_reg = 3'b111; end
            18'b101011111011011010: begin rgb_reg = 3'b111; end
            18'b101011111011100001: begin rgb_reg = 3'b111; end
            18'b101011111011100010: begin rgb_reg = 3'b111; end
            18'b101011111011100101: begin rgb_reg = 3'b111; end
            18'b101011111011100110: begin rgb_reg = 3'b111; end
            18'b101011111011101101: begin rgb_reg = 3'b111; end
            18'b101011111011101110: begin rgb_reg = 3'b111; end
            18'b101011111011111101: begin rgb_reg = 3'b111; end
            18'b101011111011111110: begin rgb_reg = 3'b111; end
            18'b101011111100000101: begin rgb_reg = 3'b111; end
            18'b101011111100000110: begin rgb_reg = 3'b111; end
            18'b101011111100001001: begin rgb_reg = 3'b111; end
            18'b101011111100001010: begin rgb_reg = 3'b111; end
            18'b101011111100001111: begin rgb_reg = 3'b111; end
            18'b101011111100010000: begin rgb_reg = 3'b111; end
            18'b101011111100010001: begin rgb_reg = 3'b111; end
            18'b101011111100010010: begin rgb_reg = 3'b111; end
            18'b101011111100010011: begin rgb_reg = 3'b111; end
            18'b101011111100010100: begin rgb_reg = 3'b111; end
            18'b101011111100010101: begin rgb_reg = 3'b111; end
            18'b101011111100010110: begin rgb_reg = 3'b111; end
            18'b101011111100011001: begin rgb_reg = 3'b111; end
            18'b101011111100011010: begin rgb_reg = 3'b111; end
            18'b101011111100100001: begin rgb_reg = 3'b111; end
            18'b101011111100100010: begin rgb_reg = 3'b111; end
            18'b101011111100100101: begin rgb_reg = 3'b111; end
            18'b101011111100100110: begin rgb_reg = 3'b111; end
            18'b101011111100101101: begin rgb_reg = 3'b111; end
            18'b101011111100101110: begin rgb_reg = 3'b111; end
            18'b101011111100111001: begin rgb_reg = 3'b111; end
            18'b101011111100111010: begin rgb_reg = 3'b111; end
            18'b101011111100111101: begin rgb_reg = 3'b111; end
            18'b101011111100111110: begin rgb_reg = 3'b111; end
            18'b101011111101000101: begin rgb_reg = 3'b111; end
            18'b101011111101000110: begin rgb_reg = 3'b111; end
            18'b101011111101001011: begin rgb_reg = 3'b111; end
            18'b101011111101001100: begin rgb_reg = 3'b111; end
            18'b101011111101010001: begin rgb_reg = 3'b111; end
            18'b101011111101010010: begin rgb_reg = 3'b111; end
            18'b101011111101011001: begin rgb_reg = 3'b111; end
            18'b101011111101011010: begin rgb_reg = 3'b111; end
            18'b101011111101011101: begin rgb_reg = 3'b111; end
            18'b101011111101011110: begin rgb_reg = 3'b111; end
            18'b101011111101100001: begin rgb_reg = 3'b111; end
            18'b101011111101100010: begin rgb_reg = 3'b111; end
            18'b101011111101101101: begin rgb_reg = 3'b111; end
            18'b101011111101101110: begin rgb_reg = 3'b111; end
            18'b101011111101110101: begin rgb_reg = 3'b111; end
            18'b101011111101110110: begin rgb_reg = 3'b111; end
            18'b101100000010001001: begin rgb_reg = 3'b111; end
            18'b101100000010001010: begin rgb_reg = 3'b111; end
            18'b101100000010010001: begin rgb_reg = 3'b111; end
            18'b101100000010010010: begin rgb_reg = 3'b111; end
            18'b101100000010010101: begin rgb_reg = 3'b111; end
            18'b101100000010010110: begin rgb_reg = 3'b111; end
            18'b101100000010011101: begin rgb_reg = 3'b111; end
            18'b101100000010011110: begin rgb_reg = 3'b111; end
            18'b101100000010100011: begin rgb_reg = 3'b111; end
            18'b101100000010100100: begin rgb_reg = 3'b111; end
            18'b101100000010101001: begin rgb_reg = 3'b111; end
            18'b101100000010101010: begin rgb_reg = 3'b111; end
            18'b101100000010110001: begin rgb_reg = 3'b111; end
            18'b101100000010110010: begin rgb_reg = 3'b111; end
            18'b101100000010110101: begin rgb_reg = 3'b111; end
            18'b101100000010110110: begin rgb_reg = 3'b111; end
            18'b101100000010111101: begin rgb_reg = 3'b111; end
            18'b101100000010111110: begin rgb_reg = 3'b111; end
            18'b101100000011000001: begin rgb_reg = 3'b111; end
            18'b101100000011000010: begin rgb_reg = 3'b111; end
            18'b101100000011000011: begin rgb_reg = 3'b111; end
            18'b101100000011000100: begin rgb_reg = 3'b111; end
            18'b101100000011000101: begin rgb_reg = 3'b111; end
            18'b101100000011000110: begin rgb_reg = 3'b111; end
            18'b101100000011000111: begin rgb_reg = 3'b111; end
            18'b101100000011001000: begin rgb_reg = 3'b111; end
            18'b101100000011001101: begin rgb_reg = 3'b111; end
            18'b101100000011001110: begin rgb_reg = 3'b111; end
            18'b101100000011010101: begin rgb_reg = 3'b111; end
            18'b101100000011010110: begin rgb_reg = 3'b111; end
            18'b101100000011011001: begin rgb_reg = 3'b111; end
            18'b101100000011011010: begin rgb_reg = 3'b111; end
            18'b101100000011100001: begin rgb_reg = 3'b111; end
            18'b101100000011100010: begin rgb_reg = 3'b111; end
            18'b101100000011100101: begin rgb_reg = 3'b111; end
            18'b101100000011100110: begin rgb_reg = 3'b111; end
            18'b101100000011101101: begin rgb_reg = 3'b111; end
            18'b101100000011101110: begin rgb_reg = 3'b111; end
            18'b101100000011111101: begin rgb_reg = 3'b111; end
            18'b101100000011111110: begin rgb_reg = 3'b111; end
            18'b101100000100000101: begin rgb_reg = 3'b111; end
            18'b101100000100000110: begin rgb_reg = 3'b111; end
            18'b101100000100001001: begin rgb_reg = 3'b111; end
            18'b101100000100001010: begin rgb_reg = 3'b111; end
            18'b101100000100001111: begin rgb_reg = 3'b111; end
            18'b101100000100010000: begin rgb_reg = 3'b111; end
            18'b101100000100010001: begin rgb_reg = 3'b111; end
            18'b101100000100010010: begin rgb_reg = 3'b111; end
            18'b101100000100010011: begin rgb_reg = 3'b111; end
            18'b101100000100010100: begin rgb_reg = 3'b111; end
            18'b101100000100010101: begin rgb_reg = 3'b111; end
            18'b101100000100010110: begin rgb_reg = 3'b111; end
            18'b101100000100011001: begin rgb_reg = 3'b111; end
            18'b101100000100011010: begin rgb_reg = 3'b111; end
            18'b101100000100100001: begin rgb_reg = 3'b111; end
            18'b101100000100100010: begin rgb_reg = 3'b111; end
            18'b101100000100100101: begin rgb_reg = 3'b111; end
            18'b101100000100100110: begin rgb_reg = 3'b111; end
            18'b101100000100101101: begin rgb_reg = 3'b111; end
            18'b101100000100101110: begin rgb_reg = 3'b111; end
            18'b101100000100111001: begin rgb_reg = 3'b111; end
            18'b101100000100111010: begin rgb_reg = 3'b111; end
            18'b101100000100111101: begin rgb_reg = 3'b111; end
            18'b101100000100111110: begin rgb_reg = 3'b111; end
            18'b101100000101000101: begin rgb_reg = 3'b111; end
            18'b101100000101000110: begin rgb_reg = 3'b111; end
            18'b101100000101001011: begin rgb_reg = 3'b111; end
            18'b101100000101001100: begin rgb_reg = 3'b111; end
            18'b101100000101010001: begin rgb_reg = 3'b111; end
            18'b101100000101010010: begin rgb_reg = 3'b111; end
            18'b101100000101011001: begin rgb_reg = 3'b111; end
            18'b101100000101011010: begin rgb_reg = 3'b111; end
            18'b101100000101011101: begin rgb_reg = 3'b111; end
            18'b101100000101011110: begin rgb_reg = 3'b111; end
            18'b101100000101100001: begin rgb_reg = 3'b111; end
            18'b101100000101100010: begin rgb_reg = 3'b111; end
            18'b101100000101101101: begin rgb_reg = 3'b111; end
            18'b101100000101101110: begin rgb_reg = 3'b111; end
            18'b101100000101110101: begin rgb_reg = 3'b111; end
            18'b101100000101110110: begin rgb_reg = 3'b111; end
            18'b101100001010001001: begin rgb_reg = 3'b111; end
            18'b101100001010001010: begin rgb_reg = 3'b111; end
            18'b101100001010010001: begin rgb_reg = 3'b111; end
            18'b101100001010010010: begin rgb_reg = 3'b111; end
            18'b101100001010010111: begin rgb_reg = 3'b111; end
            18'b101100001010011000: begin rgb_reg = 3'b111; end
            18'b101100001010011001: begin rgb_reg = 3'b111; end
            18'b101100001010011010: begin rgb_reg = 3'b111; end
            18'b101100001010011011: begin rgb_reg = 3'b111; end
            18'b101100001010011100: begin rgb_reg = 3'b111; end
            18'b101100001010011101: begin rgb_reg = 3'b111; end
            18'b101100001010011110: begin rgb_reg = 3'b111; end
            18'b101100001010100101: begin rgb_reg = 3'b111; end
            18'b101100001010100110: begin rgb_reg = 3'b111; end
            18'b101100001010101001: begin rgb_reg = 3'b111; end
            18'b101100001010101010: begin rgb_reg = 3'b111; end
            18'b101100001010110001: begin rgb_reg = 3'b111; end
            18'b101100001010110010: begin rgb_reg = 3'b111; end
            18'b101100001010110111: begin rgb_reg = 3'b111; end
            18'b101100001010111000: begin rgb_reg = 3'b111; end
            18'b101100001010111001: begin rgb_reg = 3'b111; end
            18'b101100001010111010: begin rgb_reg = 3'b111; end
            18'b101100001010111011: begin rgb_reg = 3'b111; end
            18'b101100001010111100: begin rgb_reg = 3'b111; end
            18'b101100001010111101: begin rgb_reg = 3'b111; end
            18'b101100001010111110: begin rgb_reg = 3'b111; end
            18'b101100001011000001: begin rgb_reg = 3'b111; end
            18'b101100001011000010: begin rgb_reg = 3'b111; end
            18'b101100001011001101: begin rgb_reg = 3'b111; end
            18'b101100001011001110: begin rgb_reg = 3'b111; end
            18'b101100001011010101: begin rgb_reg = 3'b111; end
            18'b101100001011010110: begin rgb_reg = 3'b111; end
            18'b101100001011011011: begin rgb_reg = 3'b111; end
            18'b101100001011011100: begin rgb_reg = 3'b111; end
            18'b101100001011011101: begin rgb_reg = 3'b111; end
            18'b101100001011011110: begin rgb_reg = 3'b111; end
            18'b101100001011011111: begin rgb_reg = 3'b111; end
            18'b101100001011100000: begin rgb_reg = 3'b111; end
            18'b101100001011100001: begin rgb_reg = 3'b111; end
            18'b101100001011100010: begin rgb_reg = 3'b111; end
            18'b101100001011100101: begin rgb_reg = 3'b111; end
            18'b101100001011100110: begin rgb_reg = 3'b111; end
            18'b101100001011101101: begin rgb_reg = 3'b111; end
            18'b101100001011101110: begin rgb_reg = 3'b111; end
            18'b101100001011111101: begin rgb_reg = 3'b111; end
            18'b101100001011111110: begin rgb_reg = 3'b111; end
            18'b101100001100000101: begin rgb_reg = 3'b111; end
            18'b101100001100000110: begin rgb_reg = 3'b111; end
            18'b101100001100001001: begin rgb_reg = 3'b111; end
            18'b101100001100001010: begin rgb_reg = 3'b111; end
            18'b101100001100010101: begin rgb_reg = 3'b111; end
            18'b101100001100010110: begin rgb_reg = 3'b111; end
            18'b101100001100011011: begin rgb_reg = 3'b111; end
            18'b101100001100011100: begin rgb_reg = 3'b111; end
            18'b101100001100011101: begin rgb_reg = 3'b111; end
            18'b101100001100011110: begin rgb_reg = 3'b111; end
            18'b101100001100011111: begin rgb_reg = 3'b111; end
            18'b101100001100100000: begin rgb_reg = 3'b111; end
            18'b101100001100100101: begin rgb_reg = 3'b111; end
            18'b101100001100100110: begin rgb_reg = 3'b111; end
            18'b101100001100101101: begin rgb_reg = 3'b111; end
            18'b101100001100101110: begin rgb_reg = 3'b111; end
            18'b101100001100110001: begin rgb_reg = 3'b111; end
            18'b101100001100110010: begin rgb_reg = 3'b111; end
            18'b101100001100110011: begin rgb_reg = 3'b111; end
            18'b101100001100110100: begin rgb_reg = 3'b111; end
            18'b101100001100110101: begin rgb_reg = 3'b111; end
            18'b101100001100110110: begin rgb_reg = 3'b111; end
            18'b101100001100110111: begin rgb_reg = 3'b111; end
            18'b101100001100111000: begin rgb_reg = 3'b111; end
            18'b101100001100111111: begin rgb_reg = 3'b111; end
            18'b101100001101000000: begin rgb_reg = 3'b111; end
            18'b101100001101000001: begin rgb_reg = 3'b111; end
            18'b101100001101000010: begin rgb_reg = 3'b111; end
            18'b101100001101000011: begin rgb_reg = 3'b111; end
            18'b101100001101000100: begin rgb_reg = 3'b111; end
            18'b101100001101000101: begin rgb_reg = 3'b111; end
            18'b101100001101000110: begin rgb_reg = 3'b111; end
            18'b101100001101001101: begin rgb_reg = 3'b111; end
            18'b101100001101001110: begin rgb_reg = 3'b111; end
            18'b101100001101010001: begin rgb_reg = 3'b111; end
            18'b101100001101010010: begin rgb_reg = 3'b111; end
            18'b101100001101011001: begin rgb_reg = 3'b111; end
            18'b101100001101011010: begin rgb_reg = 3'b111; end
            18'b101100001101011101: begin rgb_reg = 3'b111; end
            18'b101100001101011110: begin rgb_reg = 3'b111; end
            18'b101100001101100011: begin rgb_reg = 3'b111; end
            18'b101100001101100100: begin rgb_reg = 3'b111; end
            18'b101100001101100101: begin rgb_reg = 3'b111; end
            18'b101100001101100110: begin rgb_reg = 3'b111; end
            18'b101100001101100111: begin rgb_reg = 3'b111; end
            18'b101100001101101000: begin rgb_reg = 3'b111; end
            18'b101100001101101001: begin rgb_reg = 3'b111; end
            18'b101100001101101010: begin rgb_reg = 3'b111; end
            18'b101100001101101101: begin rgb_reg = 3'b111; end
            18'b101100001101101110: begin rgb_reg = 3'b111; end
            18'b101100001101110101: begin rgb_reg = 3'b111; end
            18'b101100001101110110: begin rgb_reg = 3'b111; end
            18'b101100010010001001: begin rgb_reg = 3'b111; end
            18'b101100010010001010: begin rgb_reg = 3'b111; end
            18'b101100010010010001: begin rgb_reg = 3'b111; end
            18'b101100010010010010: begin rgb_reg = 3'b111; end
            18'b101100010010010111: begin rgb_reg = 3'b111; end
            18'b101100010010011000: begin rgb_reg = 3'b111; end
            18'b101100010010011001: begin rgb_reg = 3'b111; end
            18'b101100010010011010: begin rgb_reg = 3'b111; end
            18'b101100010010011011: begin rgb_reg = 3'b111; end
            18'b101100010010011100: begin rgb_reg = 3'b111; end
            18'b101100010010011101: begin rgb_reg = 3'b111; end
            18'b101100010010011110: begin rgb_reg = 3'b111; end
            18'b101100010010100101: begin rgb_reg = 3'b111; end
            18'b101100010010100110: begin rgb_reg = 3'b111; end
            18'b101100010010101001: begin rgb_reg = 3'b111; end
            18'b101100010010101010: begin rgb_reg = 3'b111; end
            18'b101100010010110001: begin rgb_reg = 3'b111; end
            18'b101100010010110010: begin rgb_reg = 3'b111; end
            18'b101100010010110111: begin rgb_reg = 3'b111; end
            18'b101100010010111000: begin rgb_reg = 3'b111; end
            18'b101100010010111001: begin rgb_reg = 3'b111; end
            18'b101100010010111010: begin rgb_reg = 3'b111; end
            18'b101100010010111011: begin rgb_reg = 3'b111; end
            18'b101100010010111100: begin rgb_reg = 3'b111; end
            18'b101100010010111101: begin rgb_reg = 3'b111; end
            18'b101100010010111110: begin rgb_reg = 3'b111; end
            18'b101100010011000001: begin rgb_reg = 3'b111; end
            18'b101100010011000010: begin rgb_reg = 3'b111; end
            18'b101100010011001101: begin rgb_reg = 3'b111; end
            18'b101100010011001110: begin rgb_reg = 3'b111; end
            18'b101100010011010101: begin rgb_reg = 3'b111; end
            18'b101100010011010110: begin rgb_reg = 3'b111; end
            18'b101100010011011011: begin rgb_reg = 3'b111; end
            18'b101100010011011100: begin rgb_reg = 3'b111; end
            18'b101100010011011101: begin rgb_reg = 3'b111; end
            18'b101100010011011110: begin rgb_reg = 3'b111; end
            18'b101100010011011111: begin rgb_reg = 3'b111; end
            18'b101100010011100000: begin rgb_reg = 3'b111; end
            18'b101100010011100001: begin rgb_reg = 3'b111; end
            18'b101100010011100010: begin rgb_reg = 3'b111; end
            18'b101100010011100101: begin rgb_reg = 3'b111; end
            18'b101100010011100110: begin rgb_reg = 3'b111; end
            18'b101100010011101101: begin rgb_reg = 3'b111; end
            18'b101100010011101110: begin rgb_reg = 3'b111; end
            18'b101100010011111101: begin rgb_reg = 3'b111; end
            18'b101100010011111110: begin rgb_reg = 3'b111; end
            18'b101100010100000101: begin rgb_reg = 3'b111; end
            18'b101100010100000110: begin rgb_reg = 3'b111; end
            18'b101100010100001001: begin rgb_reg = 3'b111; end
            18'b101100010100001010: begin rgb_reg = 3'b111; end
            18'b101100010100010101: begin rgb_reg = 3'b111; end
            18'b101100010100010110: begin rgb_reg = 3'b111; end
            18'b101100010100011011: begin rgb_reg = 3'b111; end
            18'b101100010100011100: begin rgb_reg = 3'b111; end
            18'b101100010100011101: begin rgb_reg = 3'b111; end
            18'b101100010100011110: begin rgb_reg = 3'b111; end
            18'b101100010100011111: begin rgb_reg = 3'b111; end
            18'b101100010100100000: begin rgb_reg = 3'b111; end
            18'b101100010100100101: begin rgb_reg = 3'b111; end
            18'b101100010100100110: begin rgb_reg = 3'b111; end
            18'b101100010100101101: begin rgb_reg = 3'b111; end
            18'b101100010100101110: begin rgb_reg = 3'b111; end
            18'b101100010100110001: begin rgb_reg = 3'b111; end
            18'b101100010100110010: begin rgb_reg = 3'b111; end
            18'b101100010100110011: begin rgb_reg = 3'b111; end
            18'b101100010100110100: begin rgb_reg = 3'b111; end
            18'b101100010100110101: begin rgb_reg = 3'b111; end
            18'b101100010100110110: begin rgb_reg = 3'b111; end
            18'b101100010100110111: begin rgb_reg = 3'b111; end
            18'b101100010100111000: begin rgb_reg = 3'b111; end
            18'b101100010100111111: begin rgb_reg = 3'b111; end
            18'b101100010101000000: begin rgb_reg = 3'b111; end
            18'b101100010101000001: begin rgb_reg = 3'b111; end
            18'b101100010101000010: begin rgb_reg = 3'b111; end
            18'b101100010101000011: begin rgb_reg = 3'b111; end
            18'b101100010101000100: begin rgb_reg = 3'b111; end
            18'b101100010101000101: begin rgb_reg = 3'b111; end
            18'b101100010101000110: begin rgb_reg = 3'b111; end
            18'b101100010101001101: begin rgb_reg = 3'b111; end
            18'b101100010101001110: begin rgb_reg = 3'b111; end
            18'b101100010101010001: begin rgb_reg = 3'b111; end
            18'b101100010101010010: begin rgb_reg = 3'b111; end
            18'b101100010101011001: begin rgb_reg = 3'b111; end
            18'b101100010101011010: begin rgb_reg = 3'b111; end
            18'b101100010101011101: begin rgb_reg = 3'b111; end
            18'b101100010101011110: begin rgb_reg = 3'b111; end
            18'b101100010101100011: begin rgb_reg = 3'b111; end
            18'b101100010101100100: begin rgb_reg = 3'b111; end
            18'b101100010101100101: begin rgb_reg = 3'b111; end
            18'b101100010101100110: begin rgb_reg = 3'b111; end
            18'b101100010101100111: begin rgb_reg = 3'b111; end
            18'b101100010101101000: begin rgb_reg = 3'b111; end
            18'b101100010101101001: begin rgb_reg = 3'b111; end
            18'b101100010101101010: begin rgb_reg = 3'b111; end
            18'b101100010101101101: begin rgb_reg = 3'b111; end
            18'b101100010101101110: begin rgb_reg = 3'b111; end
            18'b101100010101110101: begin rgb_reg = 3'b111; end
            18'b101100010101110110: begin rgb_reg = 3'b111; end
            18'b101100011011000001: begin rgb_reg = 3'b111; end
            18'b101100011011000010: begin rgb_reg = 3'b111; end
            18'b101100011100001101: begin rgb_reg = 3'b111; end
            18'b101100011100001110: begin rgb_reg = 3'b111; end
            18'b101100011100001111: begin rgb_reg = 3'b111; end
            18'b101100011100010000: begin rgb_reg = 3'b111; end
            18'b101100011100010001: begin rgb_reg = 3'b111; end
            18'b101100011100010010: begin rgb_reg = 3'b111; end
            18'b101100011100010011: begin rgb_reg = 3'b111; end
            18'b101100011100010100: begin rgb_reg = 3'b111; end
            18'b101100100011000001: begin rgb_reg = 3'b111; end
            18'b101100100011000010: begin rgb_reg = 3'b111; end
            18'b101100100100001101: begin rgb_reg = 3'b111; end
            18'b101100100100001110: begin rgb_reg = 3'b111; end
            18'b101100100100001111: begin rgb_reg = 3'b111; end
            18'b101100100100010000: begin rgb_reg = 3'b111; end
            18'b101100100100010001: begin rgb_reg = 3'b111; end
            18'b101100100100010010: begin rgb_reg = 3'b111; end
            18'b101100100100010011: begin rgb_reg = 3'b111; end
            18'b101100100100010100: begin rgb_reg = 3'b111; end
            18'b101111000011000010: begin rgb_reg = 3'b111; end
            18'b101111000011000011: begin rgb_reg = 3'b111; end
            18'b101111000011000100: begin rgb_reg = 3'b111; end
            18'b101111000011000101: begin rgb_reg = 3'b111; end
            18'b101111000011000110: begin rgb_reg = 3'b111; end
            18'b101111000011001101: begin rgb_reg = 3'b111; end
            18'b101111000011001110: begin rgb_reg = 3'b111; end
            18'b101111000011001111: begin rgb_reg = 3'b111; end
            18'b101111000011010000: begin rgb_reg = 3'b111; end
            18'b101111000011010001: begin rgb_reg = 3'b111; end
            18'b101111000011010010: begin rgb_reg = 3'b111; end
            18'b101111000011010011: begin rgb_reg = 3'b111; end
            18'b101111000011011011: begin rgb_reg = 3'b111; end
            18'b101111000011011100: begin rgb_reg = 3'b111; end
            18'b101111000011011101: begin rgb_reg = 3'b111; end
            18'b101111000011011110: begin rgb_reg = 3'b111; end
            18'b101111000011011111: begin rgb_reg = 3'b111; end
            18'b101111000011100000: begin rgb_reg = 3'b111; end
            18'b101111000011100001: begin rgb_reg = 3'b111; end
            18'b101111000011101000: begin rgb_reg = 3'b111; end
            18'b101111000011101001: begin rgb_reg = 3'b111; end
            18'b101111000011101010: begin rgb_reg = 3'b111; end
            18'b101111000011101011: begin rgb_reg = 3'b111; end
            18'b101111000011101100: begin rgb_reg = 3'b111; end
            18'b101111000011101101: begin rgb_reg = 3'b111; end
            18'b101111000011101110: begin rgb_reg = 3'b111; end
            18'b101111000011110110: begin rgb_reg = 3'b111; end
            18'b101111000011110111: begin rgb_reg = 3'b111; end
            18'b101111000011111000: begin rgb_reg = 3'b111; end
            18'b101111000011111001: begin rgb_reg = 3'b111; end
            18'b101111000011111010: begin rgb_reg = 3'b111; end
            18'b101111000011111011: begin rgb_reg = 3'b111; end
            18'b101111000011111100: begin rgb_reg = 3'b111; end
            18'b101111000100000011: begin rgb_reg = 3'b111; end
            18'b101111000100000100: begin rgb_reg = 3'b111; end
            18'b101111000100000101: begin rgb_reg = 3'b111; end
            18'b101111000100000110: begin rgb_reg = 3'b111; end
            18'b101111000100000111: begin rgb_reg = 3'b111; end
            18'b101111000100001000: begin rgb_reg = 3'b111; end
            18'b101111000100001001: begin rgb_reg = 3'b111; end
            18'b101111000100010001: begin rgb_reg = 3'b111; end
            18'b101111000100010010: begin rgb_reg = 3'b111; end
            18'b101111000100010011: begin rgb_reg = 3'b111; end
            18'b101111000100010100: begin rgb_reg = 3'b111; end
            18'b101111000100010101: begin rgb_reg = 3'b111; end
            18'b101111000100010110: begin rgb_reg = 3'b111; end
            18'b101111000100010111: begin rgb_reg = 3'b111; end
            18'b101111000100100011: begin rgb_reg = 3'b111; end
            18'b101111000100100100: begin rgb_reg = 3'b111; end
            18'b101111000100100101: begin rgb_reg = 3'b111; end
            18'b101111000100100110: begin rgb_reg = 3'b111; end
            18'b101111000100100111: begin rgb_reg = 3'b111; end
            18'b101111000100101100: begin rgb_reg = 3'b111; end
            18'b101111000100101101: begin rgb_reg = 3'b111; end
            18'b101111000100101110: begin rgb_reg = 3'b111; end
            18'b101111000100101111: begin rgb_reg = 3'b111; end
            18'b101111000100110000: begin rgb_reg = 3'b111; end
            18'b101111000100110001: begin rgb_reg = 3'b111; end
            18'b101111000100110010: begin rgb_reg = 3'b111; end
            18'b101111000100111100: begin rgb_reg = 3'b111; end
            18'b101111000100111101: begin rgb_reg = 3'b111; end
            18'b101111001011000010: begin rgb_reg = 3'b111; end
            18'b101111001011000011: begin rgb_reg = 3'b111; end
            18'b101111001011000100: begin rgb_reg = 3'b111; end
            18'b101111001011000101: begin rgb_reg = 3'b111; end
            18'b101111001011000110: begin rgb_reg = 3'b111; end
            18'b101111001011001101: begin rgb_reg = 3'b111; end
            18'b101111001011001110: begin rgb_reg = 3'b111; end
            18'b101111001011001111: begin rgb_reg = 3'b111; end
            18'b101111001011010000: begin rgb_reg = 3'b111; end
            18'b101111001011010001: begin rgb_reg = 3'b111; end
            18'b101111001011010010: begin rgb_reg = 3'b111; end
            18'b101111001011010011: begin rgb_reg = 3'b111; end
            18'b101111001011011011: begin rgb_reg = 3'b111; end
            18'b101111001011011100: begin rgb_reg = 3'b111; end
            18'b101111001011011101: begin rgb_reg = 3'b111; end
            18'b101111001011011110: begin rgb_reg = 3'b111; end
            18'b101111001011011111: begin rgb_reg = 3'b111; end
            18'b101111001011100000: begin rgb_reg = 3'b111; end
            18'b101111001011100001: begin rgb_reg = 3'b111; end
            18'b101111001011101000: begin rgb_reg = 3'b111; end
            18'b101111001011101001: begin rgb_reg = 3'b111; end
            18'b101111001011101010: begin rgb_reg = 3'b111; end
            18'b101111001011101011: begin rgb_reg = 3'b111; end
            18'b101111001011101100: begin rgb_reg = 3'b111; end
            18'b101111001011101101: begin rgb_reg = 3'b111; end
            18'b101111001011101110: begin rgb_reg = 3'b111; end
            18'b101111001011110110: begin rgb_reg = 3'b111; end
            18'b101111001011110111: begin rgb_reg = 3'b111; end
            18'b101111001011111000: begin rgb_reg = 3'b111; end
            18'b101111001011111001: begin rgb_reg = 3'b111; end
            18'b101111001011111010: begin rgb_reg = 3'b111; end
            18'b101111001011111011: begin rgb_reg = 3'b111; end
            18'b101111001011111100: begin rgb_reg = 3'b111; end
            18'b101111001100000011: begin rgb_reg = 3'b111; end
            18'b101111001100000100: begin rgb_reg = 3'b111; end
            18'b101111001100000101: begin rgb_reg = 3'b111; end
            18'b101111001100000110: begin rgb_reg = 3'b111; end
            18'b101111001100000111: begin rgb_reg = 3'b111; end
            18'b101111001100001000: begin rgb_reg = 3'b111; end
            18'b101111001100001001: begin rgb_reg = 3'b111; end
            18'b101111001100010001: begin rgb_reg = 3'b111; end
            18'b101111001100010010: begin rgb_reg = 3'b111; end
            18'b101111001100010011: begin rgb_reg = 3'b111; end
            18'b101111001100010100: begin rgb_reg = 3'b111; end
            18'b101111001100010101: begin rgb_reg = 3'b111; end
            18'b101111001100010110: begin rgb_reg = 3'b111; end
            18'b101111001100010111: begin rgb_reg = 3'b111; end
            18'b101111001100100011: begin rgb_reg = 3'b111; end
            18'b101111001100100100: begin rgb_reg = 3'b111; end
            18'b101111001100100101: begin rgb_reg = 3'b111; end
            18'b101111001100100110: begin rgb_reg = 3'b111; end
            18'b101111001100100111: begin rgb_reg = 3'b111; end
            18'b101111001100101100: begin rgb_reg = 3'b111; end
            18'b101111001100101101: begin rgb_reg = 3'b111; end
            18'b101111001100101110: begin rgb_reg = 3'b111; end
            18'b101111001100101111: begin rgb_reg = 3'b111; end
            18'b101111001100110000: begin rgb_reg = 3'b111; end
            18'b101111001100110001: begin rgb_reg = 3'b111; end
            18'b101111001100110010: begin rgb_reg = 3'b111; end
            18'b101111001100111100: begin rgb_reg = 3'b111; end
            18'b101111001100111101: begin rgb_reg = 3'b111; end
            18'b101111010011000000: begin rgb_reg = 3'b111; end
            18'b101111010011000001: begin rgb_reg = 3'b111; end
            18'b101111010011001011: begin rgb_reg = 3'b111; end
            18'b101111010011001100: begin rgb_reg = 3'b111; end
            18'b101111010011001101: begin rgb_reg = 3'b111; end
            18'b101111010011010100: begin rgb_reg = 3'b111; end
            18'b101111010011010101: begin rgb_reg = 3'b111; end
            18'b101111010011011001: begin rgb_reg = 3'b111; end
            18'b101111010011011010: begin rgb_reg = 3'b111; end
            18'b101111010011100010: begin rgb_reg = 3'b111; end
            18'b101111010011100011: begin rgb_reg = 3'b111; end
            18'b101111010011100110: begin rgb_reg = 3'b111; end
            18'b101111010011100111: begin rgb_reg = 3'b111; end
            18'b101111010011101000: begin rgb_reg = 3'b111; end
            18'b101111010011101111: begin rgb_reg = 3'b111; end
            18'b101111010011110000: begin rgb_reg = 3'b111; end
            18'b101111010011110100: begin rgb_reg = 3'b111; end
            18'b101111010011110101: begin rgb_reg = 3'b111; end
            18'b101111010011111101: begin rgb_reg = 3'b111; end
            18'b101111010011111110: begin rgb_reg = 3'b111; end
            18'b101111010100000001: begin rgb_reg = 3'b111; end
            18'b101111010100000010: begin rgb_reg = 3'b111; end
            18'b101111010100000011: begin rgb_reg = 3'b111; end
            18'b101111010100001010: begin rgb_reg = 3'b111; end
            18'b101111010100001011: begin rgb_reg = 3'b111; end
            18'b101111010100001111: begin rgb_reg = 3'b111; end
            18'b101111010100010000: begin rgb_reg = 3'b111; end
            18'b101111010100011000: begin rgb_reg = 3'b111; end
            18'b101111010100011001: begin rgb_reg = 3'b111; end
            18'b101111010100100001: begin rgb_reg = 3'b111; end
            18'b101111010100100010: begin rgb_reg = 3'b111; end
            18'b101111010100100101: begin rgb_reg = 3'b111; end
            18'b101111010100100110: begin rgb_reg = 3'b111; end
            18'b101111010100100111: begin rgb_reg = 3'b111; end
            18'b101111010100101010: begin rgb_reg = 3'b111; end
            18'b101111010100101011: begin rgb_reg = 3'b111; end
            18'b101111010100110011: begin rgb_reg = 3'b111; end
            18'b101111010100110100: begin rgb_reg = 3'b111; end
            18'b101111010100111010: begin rgb_reg = 3'b111; end
            18'b101111010100111011: begin rgb_reg = 3'b111; end
            18'b101111010100111100: begin rgb_reg = 3'b111; end
            18'b101111010100111101: begin rgb_reg = 3'b111; end
            18'b101111011011000000: begin rgb_reg = 3'b111; end
            18'b101111011011000001: begin rgb_reg = 3'b111; end
            18'b101111011011001011: begin rgb_reg = 3'b111; end
            18'b101111011011001100: begin rgb_reg = 3'b111; end
            18'b101111011011001101: begin rgb_reg = 3'b111; end
            18'b101111011011010100: begin rgb_reg = 3'b111; end
            18'b101111011011010101: begin rgb_reg = 3'b111; end
            18'b101111011011010110: begin rgb_reg = 3'b111; end
            18'b101111011011011001: begin rgb_reg = 3'b111; end
            18'b101111011011011010: begin rgb_reg = 3'b111; end
            18'b101111011011100010: begin rgb_reg = 3'b111; end
            18'b101111011011100011: begin rgb_reg = 3'b111; end
            18'b101111011011100110: begin rgb_reg = 3'b111; end
            18'b101111011011100111: begin rgb_reg = 3'b111; end
            18'b101111011011101000: begin rgb_reg = 3'b111; end
            18'b101111011011101111: begin rgb_reg = 3'b111; end
            18'b101111011011110000: begin rgb_reg = 3'b111; end
            18'b101111011011110001: begin rgb_reg = 3'b111; end
            18'b101111011011110100: begin rgb_reg = 3'b111; end
            18'b101111011011110101: begin rgb_reg = 3'b111; end
            18'b101111011011111101: begin rgb_reg = 3'b111; end
            18'b101111011011111110: begin rgb_reg = 3'b111; end
            18'b101111011100000001: begin rgb_reg = 3'b111; end
            18'b101111011100000010: begin rgb_reg = 3'b111; end
            18'b101111011100000011: begin rgb_reg = 3'b111; end
            18'b101111011100001010: begin rgb_reg = 3'b111; end
            18'b101111011100001011: begin rgb_reg = 3'b111; end
            18'b101111011100001100: begin rgb_reg = 3'b111; end
            18'b101111011100001111: begin rgb_reg = 3'b111; end
            18'b101111011100010000: begin rgb_reg = 3'b111; end
            18'b101111011100011000: begin rgb_reg = 3'b111; end
            18'b101111011100011001: begin rgb_reg = 3'b111; end
            18'b101111011100100001: begin rgb_reg = 3'b111; end
            18'b101111011100100010: begin rgb_reg = 3'b111; end
            18'b101111011100100101: begin rgb_reg = 3'b111; end
            18'b101111011100100110: begin rgb_reg = 3'b111; end
            18'b101111011100100111: begin rgb_reg = 3'b111; end
            18'b101111011100101010: begin rgb_reg = 3'b111; end
            18'b101111011100101011: begin rgb_reg = 3'b111; end
            18'b101111011100110011: begin rgb_reg = 3'b111; end
            18'b101111011100110100: begin rgb_reg = 3'b111; end
            18'b101111011100111001: begin rgb_reg = 3'b111; end
            18'b101111011100111010: begin rgb_reg = 3'b111; end
            18'b101111011100111011: begin rgb_reg = 3'b111; end
            18'b101111011100111100: begin rgb_reg = 3'b111; end
            18'b101111011100111101: begin rgb_reg = 3'b111; end
            18'b101111100010111110: begin rgb_reg = 3'b111; end
            18'b101111100010111111: begin rgb_reg = 3'b111; end
            18'b101111100011000000: begin rgb_reg = 3'b111; end
            18'b101111100011000001: begin rgb_reg = 3'b111; end
            18'b101111100011001011: begin rgb_reg = 3'b111; end
            18'b101111100011001100: begin rgb_reg = 3'b111; end
            18'b101111100011001101: begin rgb_reg = 3'b111; end
            18'b101111100011010010: begin rgb_reg = 3'b111; end
            18'b101111100011010011: begin rgb_reg = 3'b111; end
            18'b101111100011010100: begin rgb_reg = 3'b111; end
            18'b101111100011010101: begin rgb_reg = 3'b111; end
            18'b101111100011010110: begin rgb_reg = 3'b111; end
            18'b101111100011011001: begin rgb_reg = 3'b111; end
            18'b101111100011011010: begin rgb_reg = 3'b111; end
            18'b101111100011100010: begin rgb_reg = 3'b111; end
            18'b101111100011100011: begin rgb_reg = 3'b111; end
            18'b101111100011100110: begin rgb_reg = 3'b111; end
            18'b101111100011100111: begin rgb_reg = 3'b111; end
            18'b101111100011101000: begin rgb_reg = 3'b111; end
            18'b101111100011101101: begin rgb_reg = 3'b111; end
            18'b101111100011101110: begin rgb_reg = 3'b111; end
            18'b101111100011101111: begin rgb_reg = 3'b111; end
            18'b101111100011110000: begin rgb_reg = 3'b111; end
            18'b101111100011110001: begin rgb_reg = 3'b111; end
            18'b101111100011110100: begin rgb_reg = 3'b111; end
            18'b101111100011110101: begin rgb_reg = 3'b111; end
            18'b101111100011111101: begin rgb_reg = 3'b111; end
            18'b101111100011111110: begin rgb_reg = 3'b111; end
            18'b101111100100000010: begin rgb_reg = 3'b111; end
            18'b101111100100001010: begin rgb_reg = 3'b111; end
            18'b101111100100001011: begin rgb_reg = 3'b111; end
            18'b101111100100001100: begin rgb_reg = 3'b111; end
            18'b101111100100001111: begin rgb_reg = 3'b111; end
            18'b101111100100010000: begin rgb_reg = 3'b111; end
            18'b101111100100010110: begin rgb_reg = 3'b111; end
            18'b101111100100010111: begin rgb_reg = 3'b111; end
            18'b101111100100011000: begin rgb_reg = 3'b111; end
            18'b101111100100011001: begin rgb_reg = 3'b111; end
            18'b101111100100011111: begin rgb_reg = 3'b111; end
            18'b101111100100100000: begin rgb_reg = 3'b111; end
            18'b101111100100100001: begin rgb_reg = 3'b111; end
            18'b101111100100100010: begin rgb_reg = 3'b111; end
            18'b101111100100100101: begin rgb_reg = 3'b111; end
            18'b101111100100100110: begin rgb_reg = 3'b111; end
            18'b101111100100100111: begin rgb_reg = 3'b111; end
            18'b101111100100101010: begin rgb_reg = 3'b111; end
            18'b101111100100101011: begin rgb_reg = 3'b111; end
            18'b101111100100110011: begin rgb_reg = 3'b111; end
            18'b101111100100110100: begin rgb_reg = 3'b111; end
            18'b101111100100111010: begin rgb_reg = 3'b111; end
            18'b101111100100111011: begin rgb_reg = 3'b111; end
            18'b101111100100111100: begin rgb_reg = 3'b111; end
            18'b101111100100111101: begin rgb_reg = 3'b111; end
            18'b101111101010111110: begin rgb_reg = 3'b111; end
            18'b101111101010111111: begin rgb_reg = 3'b111; end
            18'b101111101011001011: begin rgb_reg = 3'b111; end
            18'b101111101011001100: begin rgb_reg = 3'b111; end
            18'b101111101011001101: begin rgb_reg = 3'b111; end
            18'b101111101011010010: begin rgb_reg = 3'b111; end
            18'b101111101011010011: begin rgb_reg = 3'b111; end
            18'b101111101011010100: begin rgb_reg = 3'b111; end
            18'b101111101011010101: begin rgb_reg = 3'b111; end
            18'b101111101011010110: begin rgb_reg = 3'b111; end
            18'b101111101011100010: begin rgb_reg = 3'b111; end
            18'b101111101011100011: begin rgb_reg = 3'b111; end
            18'b101111101011100110: begin rgb_reg = 3'b111; end
            18'b101111101011100111: begin rgb_reg = 3'b111; end
            18'b101111101011101000: begin rgb_reg = 3'b111; end
            18'b101111101011101101: begin rgb_reg = 3'b111; end
            18'b101111101011101110: begin rgb_reg = 3'b111; end
            18'b101111101011101111: begin rgb_reg = 3'b111; end
            18'b101111101011110000: begin rgb_reg = 3'b111; end
            18'b101111101011110001: begin rgb_reg = 3'b111; end
            18'b101111101011111101: begin rgb_reg = 3'b111; end
            18'b101111101011111110: begin rgb_reg = 3'b111; end
            18'b101111101100001010: begin rgb_reg = 3'b111; end
            18'b101111101100001011: begin rgb_reg = 3'b111; end
            18'b101111101100001100: begin rgb_reg = 3'b111; end
            18'b101111101100001111: begin rgb_reg = 3'b111; end
            18'b101111101100010000: begin rgb_reg = 3'b111; end
            18'b101111101100010101: begin rgb_reg = 3'b111; end
            18'b101111101100010110: begin rgb_reg = 3'b111; end
            18'b101111101100010111: begin rgb_reg = 3'b111; end
            18'b101111101100011000: begin rgb_reg = 3'b111; end
            18'b101111101100011001: begin rgb_reg = 3'b111; end
            18'b101111101100011110: begin rgb_reg = 3'b111; end
            18'b101111101100011111: begin rgb_reg = 3'b111; end
            18'b101111101100100000: begin rgb_reg = 3'b111; end
            18'b101111101100100101: begin rgb_reg = 3'b111; end
            18'b101111101100100110: begin rgb_reg = 3'b111; end
            18'b101111101100100111: begin rgb_reg = 3'b111; end
            18'b101111101100110011: begin rgb_reg = 3'b111; end
            18'b101111101100110100: begin rgb_reg = 3'b111; end
            18'b101111101100111100: begin rgb_reg = 3'b111; end
            18'b101111101100111101: begin rgb_reg = 3'b111; end
            18'b101111110010111110: begin rgb_reg = 3'b111; end
            18'b101111110010111111: begin rgb_reg = 3'b111; end
            18'b101111110011001011: begin rgb_reg = 3'b111; end
            18'b101111110011001100: begin rgb_reg = 3'b111; end
            18'b101111110011001101: begin rgb_reg = 3'b111; end
            18'b101111110011010010: begin rgb_reg = 3'b111; end
            18'b101111110011010011: begin rgb_reg = 3'b111; end
            18'b101111110011010100: begin rgb_reg = 3'b111; end
            18'b101111110011010101: begin rgb_reg = 3'b111; end
            18'b101111110011010110: begin rgb_reg = 3'b111; end
            18'b101111110011100010: begin rgb_reg = 3'b111; end
            18'b101111110011100011: begin rgb_reg = 3'b111; end
            18'b101111110011100110: begin rgb_reg = 3'b111; end
            18'b101111110011100111: begin rgb_reg = 3'b111; end
            18'b101111110011101000: begin rgb_reg = 3'b111; end
            18'b101111110011101101: begin rgb_reg = 3'b111; end
            18'b101111110011101110: begin rgb_reg = 3'b111; end
            18'b101111110011101111: begin rgb_reg = 3'b111; end
            18'b101111110011110000: begin rgb_reg = 3'b111; end
            18'b101111110011110001: begin rgb_reg = 3'b111; end
            18'b101111110011111101: begin rgb_reg = 3'b111; end
            18'b101111110011111110: begin rgb_reg = 3'b111; end
            18'b101111110100001010: begin rgb_reg = 3'b111; end
            18'b101111110100001011: begin rgb_reg = 3'b111; end
            18'b101111110100001111: begin rgb_reg = 3'b111; end
            18'b101111110100010000: begin rgb_reg = 3'b111; end
            18'b101111110100010101: begin rgb_reg = 3'b111; end
            18'b101111110100010110: begin rgb_reg = 3'b111; end
            18'b101111110100010111: begin rgb_reg = 3'b111; end
            18'b101111110100011000: begin rgb_reg = 3'b111; end
            18'b101111110100011001: begin rgb_reg = 3'b111; end
            18'b101111110100011110: begin rgb_reg = 3'b111; end
            18'b101111110100011111: begin rgb_reg = 3'b111; end
            18'b101111110100100000: begin rgb_reg = 3'b111; end
            18'b101111110100100101: begin rgb_reg = 3'b111; end
            18'b101111110100100110: begin rgb_reg = 3'b111; end
            18'b101111110100100111: begin rgb_reg = 3'b111; end
            18'b101111110100110011: begin rgb_reg = 3'b111; end
            18'b101111110100110100: begin rgb_reg = 3'b111; end
            18'b101111110100111100: begin rgb_reg = 3'b111; end
            18'b101111110100111101: begin rgb_reg = 3'b111; end
            18'b101111111010111110: begin rgb_reg = 3'b111; end
            18'b101111111010111111: begin rgb_reg = 3'b111; end
            18'b101111111011000000: begin rgb_reg = 3'b111; end
            18'b101111111011000001: begin rgb_reg = 3'b111; end
            18'b101111111011000010: begin rgb_reg = 3'b111; end
            18'b101111111011000011: begin rgb_reg = 3'b111; end
            18'b101111111011000100: begin rgb_reg = 3'b111; end
            18'b101111111011000101: begin rgb_reg = 3'b111; end
            18'b101111111011000110: begin rgb_reg = 3'b111; end
            18'b101111111011001011: begin rgb_reg = 3'b111; end
            18'b101111111011001100: begin rgb_reg = 3'b111; end
            18'b101111111011001101: begin rgb_reg = 3'b111; end
            18'b101111111011010000: begin rgb_reg = 3'b111; end
            18'b101111111011010001: begin rgb_reg = 3'b111; end
            18'b101111111011010100: begin rgb_reg = 3'b111; end
            18'b101111111011010101: begin rgb_reg = 3'b111; end
            18'b101111111011010110: begin rgb_reg = 3'b111; end
            18'b101111111011011101: begin rgb_reg = 3'b111; end
            18'b101111111011011110: begin rgb_reg = 3'b111; end
            18'b101111111011011111: begin rgb_reg = 3'b111; end
            18'b101111111011100000: begin rgb_reg = 3'b111; end
            18'b101111111011100001: begin rgb_reg = 3'b111; end
            18'b101111111011100110: begin rgb_reg = 3'b111; end
            18'b101111111011100111: begin rgb_reg = 3'b111; end
            18'b101111111011101000: begin rgb_reg = 3'b111; end
            18'b101111111011101011: begin rgb_reg = 3'b111; end
            18'b101111111011101100: begin rgb_reg = 3'b111; end
            18'b101111111011101111: begin rgb_reg = 3'b111; end
            18'b101111111011110000: begin rgb_reg = 3'b111; end
            18'b101111111011110001: begin rgb_reg = 3'b111; end
            18'b101111111011111000: begin rgb_reg = 3'b111; end
            18'b101111111011111001: begin rgb_reg = 3'b111; end
            18'b101111111011111010: begin rgb_reg = 3'b111; end
            18'b101111111011111011: begin rgb_reg = 3'b111; end
            18'b101111111011111100: begin rgb_reg = 3'b111; end
            18'b101111111100000110: begin rgb_reg = 3'b111; end
            18'b101111111100000111: begin rgb_reg = 3'b111; end
            18'b101111111100001000: begin rgb_reg = 3'b111; end
            18'b101111111100001001: begin rgb_reg = 3'b111; end
            18'b101111111100001111: begin rgb_reg = 3'b111; end
            18'b101111111100010000: begin rgb_reg = 3'b111; end
            18'b101111111100010011: begin rgb_reg = 3'b111; end
            18'b101111111100010100: begin rgb_reg = 3'b111; end
            18'b101111111100010101: begin rgb_reg = 3'b111; end
            18'b101111111100011000: begin rgb_reg = 3'b111; end
            18'b101111111100011001: begin rgb_reg = 3'b111; end
            18'b101111111100011100: begin rgb_reg = 3'b111; end
            18'b101111111100011101: begin rgb_reg = 3'b111; end
            18'b101111111100011110: begin rgb_reg = 3'b111; end
            18'b101111111100100101: begin rgb_reg = 3'b111; end
            18'b101111111100100110: begin rgb_reg = 3'b111; end
            18'b101111111100100111: begin rgb_reg = 3'b111; end
            18'b101111111100101110: begin rgb_reg = 3'b111; end
            18'b101111111100101111: begin rgb_reg = 3'b111; end
            18'b101111111100110000: begin rgb_reg = 3'b111; end
            18'b101111111100110001: begin rgb_reg = 3'b111; end
            18'b101111111100110010: begin rgb_reg = 3'b111; end
            18'b101111111100111100: begin rgb_reg = 3'b111; end
            18'b101111111100111101: begin rgb_reg = 3'b111; end
            18'b110000000010111110: begin rgb_reg = 3'b111; end
            18'b110000000010111111: begin rgb_reg = 3'b111; end
            18'b110000000011000000: begin rgb_reg = 3'b111; end
            18'b110000000011000001: begin rgb_reg = 3'b111; end
            18'b110000000011000010: begin rgb_reg = 3'b111; end
            18'b110000000011000011: begin rgb_reg = 3'b111; end
            18'b110000000011000100: begin rgb_reg = 3'b111; end
            18'b110000000011000101: begin rgb_reg = 3'b111; end
            18'b110000000011000110: begin rgb_reg = 3'b111; end
            18'b110000000011001011: begin rgb_reg = 3'b111; end
            18'b110000000011001100: begin rgb_reg = 3'b111; end
            18'b110000000011001101: begin rgb_reg = 3'b111; end
            18'b110000000011010000: begin rgb_reg = 3'b111; end
            18'b110000000011010001: begin rgb_reg = 3'b111; end
            18'b110000000011010100: begin rgb_reg = 3'b111; end
            18'b110000000011010101: begin rgb_reg = 3'b111; end
            18'b110000000011010110: begin rgb_reg = 3'b111; end
            18'b110000000011011101: begin rgb_reg = 3'b111; end
            18'b110000000011011110: begin rgb_reg = 3'b111; end
            18'b110000000011011111: begin rgb_reg = 3'b111; end
            18'b110000000011100000: begin rgb_reg = 3'b111; end
            18'b110000000011100001: begin rgb_reg = 3'b111; end
            18'b110000000011100110: begin rgb_reg = 3'b111; end
            18'b110000000011100111: begin rgb_reg = 3'b111; end
            18'b110000000011101000: begin rgb_reg = 3'b111; end
            18'b110000000011101011: begin rgb_reg = 3'b111; end
            18'b110000000011101100: begin rgb_reg = 3'b111; end
            18'b110000000011101111: begin rgb_reg = 3'b111; end
            18'b110000000011110000: begin rgb_reg = 3'b111; end
            18'b110000000011110001: begin rgb_reg = 3'b111; end
            18'b110000000011111000: begin rgb_reg = 3'b111; end
            18'b110000000011111001: begin rgb_reg = 3'b111; end
            18'b110000000011111010: begin rgb_reg = 3'b111; end
            18'b110000000011111011: begin rgb_reg = 3'b111; end
            18'b110000000011111100: begin rgb_reg = 3'b111; end
            18'b110000000100000110: begin rgb_reg = 3'b111; end
            18'b110000000100000111: begin rgb_reg = 3'b111; end
            18'b110000000100001000: begin rgb_reg = 3'b111; end
            18'b110000000100001001: begin rgb_reg = 3'b111; end
            18'b110000000100001111: begin rgb_reg = 3'b111; end
            18'b110000000100010000: begin rgb_reg = 3'b111; end
            18'b110000000100010011: begin rgb_reg = 3'b111; end
            18'b110000000100010100: begin rgb_reg = 3'b111; end
            18'b110000000100010101: begin rgb_reg = 3'b111; end
            18'b110000000100011000: begin rgb_reg = 3'b111; end
            18'b110000000100011001: begin rgb_reg = 3'b111; end
            18'b110000000100011100: begin rgb_reg = 3'b111; end
            18'b110000000100011101: begin rgb_reg = 3'b111; end
            18'b110000000100011110: begin rgb_reg = 3'b111; end
            18'b110000000100100101: begin rgb_reg = 3'b111; end
            18'b110000000100100110: begin rgb_reg = 3'b111; end
            18'b110000000100100111: begin rgb_reg = 3'b111; end
            18'b110000000100101110: begin rgb_reg = 3'b111; end
            18'b110000000100101111: begin rgb_reg = 3'b111; end
            18'b110000000100110000: begin rgb_reg = 3'b111; end
            18'b110000000100110001: begin rgb_reg = 3'b111; end
            18'b110000000100110010: begin rgb_reg = 3'b111; end
            18'b110000000100111100: begin rgb_reg = 3'b111; end
            18'b110000000100111101: begin rgb_reg = 3'b111; end
            18'b110000001010111110: begin rgb_reg = 3'b111; end
            18'b110000001010111111: begin rgb_reg = 3'b111; end
            18'b110000001011000111: begin rgb_reg = 3'b111; end
            18'b110000001011001000: begin rgb_reg = 3'b111; end
            18'b110000001011001011: begin rgb_reg = 3'b111; end
            18'b110000001011001100: begin rgb_reg = 3'b111; end
            18'b110000001011001101: begin rgb_reg = 3'b111; end
            18'b110000001011001110: begin rgb_reg = 3'b111; end
            18'b110000001011001111: begin rgb_reg = 3'b111; end
            18'b110000001011010100: begin rgb_reg = 3'b111; end
            18'b110000001011010101: begin rgb_reg = 3'b111; end
            18'b110000001011010110: begin rgb_reg = 3'b111; end
            18'b110000001011100010: begin rgb_reg = 3'b111; end
            18'b110000001011100011: begin rgb_reg = 3'b111; end
            18'b110000001011100110: begin rgb_reg = 3'b111; end
            18'b110000001011100111: begin rgb_reg = 3'b111; end
            18'b110000001011101000: begin rgb_reg = 3'b111; end
            18'b110000001011101001: begin rgb_reg = 3'b111; end
            18'b110000001011101010: begin rgb_reg = 3'b111; end
            18'b110000001011101111: begin rgb_reg = 3'b111; end
            18'b110000001011110000: begin rgb_reg = 3'b111; end
            18'b110000001011110001: begin rgb_reg = 3'b111; end
            18'b110000001011111101: begin rgb_reg = 3'b111; end
            18'b110000001011111110: begin rgb_reg = 3'b111; end
            18'b110000001100000011: begin rgb_reg = 3'b111; end
            18'b110000001100000100: begin rgb_reg = 3'b111; end
            18'b110000001100000101: begin rgb_reg = 3'b111; end
            18'b110000001100001111: begin rgb_reg = 3'b111; end
            18'b110000001100010000: begin rgb_reg = 3'b111; end
            18'b110000001100010001: begin rgb_reg = 3'b111; end
            18'b110000001100010010: begin rgb_reg = 3'b111; end
            18'b110000001100011000: begin rgb_reg = 3'b111; end
            18'b110000001100011001: begin rgb_reg = 3'b111; end
            18'b110000001100011100: begin rgb_reg = 3'b111; end
            18'b110000001100011101: begin rgb_reg = 3'b111; end
            18'b110000001100011110: begin rgb_reg = 3'b111; end
            18'b110000001100011111: begin rgb_reg = 3'b111; end
            18'b110000001100100000: begin rgb_reg = 3'b111; end
            18'b110000001100100001: begin rgb_reg = 3'b111; end
            18'b110000001100100010: begin rgb_reg = 3'b111; end
            18'b110000001100100011: begin rgb_reg = 3'b111; end
            18'b110000001100100100: begin rgb_reg = 3'b111; end
            18'b110000001100100101: begin rgb_reg = 3'b111; end
            18'b110000001100100110: begin rgb_reg = 3'b111; end
            18'b110000001100100111: begin rgb_reg = 3'b111; end
            18'b110000001100101100: begin rgb_reg = 3'b111; end
            18'b110000001100101101: begin rgb_reg = 3'b111; end
            18'b110000001100111100: begin rgb_reg = 3'b111; end
            18'b110000001100111101: begin rgb_reg = 3'b111; end
            18'b110000010010111110: begin rgb_reg = 3'b111; end
            18'b110000010010111111: begin rgb_reg = 3'b111; end
            18'b110000010011000111: begin rgb_reg = 3'b111; end
            18'b110000010011001000: begin rgb_reg = 3'b111; end
            18'b110000010011001011: begin rgb_reg = 3'b111; end
            18'b110000010011001100: begin rgb_reg = 3'b111; end
            18'b110000010011001101: begin rgb_reg = 3'b111; end
            18'b110000010011001110: begin rgb_reg = 3'b111; end
            18'b110000010011001111: begin rgb_reg = 3'b111; end
            18'b110000010011010100: begin rgb_reg = 3'b111; end
            18'b110000010011010101: begin rgb_reg = 3'b111; end
            18'b110000010011010110: begin rgb_reg = 3'b111; end
            18'b110000010011100010: begin rgb_reg = 3'b111; end
            18'b110000010011100011: begin rgb_reg = 3'b111; end
            18'b110000010011100110: begin rgb_reg = 3'b111; end
            18'b110000010011100111: begin rgb_reg = 3'b111; end
            18'b110000010011101000: begin rgb_reg = 3'b111; end
            18'b110000010011101001: begin rgb_reg = 3'b111; end
            18'b110000010011101010: begin rgb_reg = 3'b111; end
            18'b110000010011101111: begin rgb_reg = 3'b111; end
            18'b110000010011110000: begin rgb_reg = 3'b111; end
            18'b110000010011110001: begin rgb_reg = 3'b111; end
            18'b110000010011111101: begin rgb_reg = 3'b111; end
            18'b110000010011111110: begin rgb_reg = 3'b111; end
            18'b110000010100000011: begin rgb_reg = 3'b111; end
            18'b110000010100000100: begin rgb_reg = 3'b111; end
            18'b110000010100000101: begin rgb_reg = 3'b111; end
            18'b110000010100001111: begin rgb_reg = 3'b111; end
            18'b110000010100010000: begin rgb_reg = 3'b111; end
            18'b110000010100010001: begin rgb_reg = 3'b111; end
            18'b110000010100010010: begin rgb_reg = 3'b111; end
            18'b110000010100011000: begin rgb_reg = 3'b111; end
            18'b110000010100011001: begin rgb_reg = 3'b111; end
            18'b110000010100011100: begin rgb_reg = 3'b111; end
            18'b110000010100011101: begin rgb_reg = 3'b111; end
            18'b110000010100011110: begin rgb_reg = 3'b111; end
            18'b110000010100011111: begin rgb_reg = 3'b111; end
            18'b110000010100100000: begin rgb_reg = 3'b111; end
            18'b110000010100100001: begin rgb_reg = 3'b111; end
            18'b110000010100100010: begin rgb_reg = 3'b111; end
            18'b110000010100100011: begin rgb_reg = 3'b111; end
            18'b110000010100100100: begin rgb_reg = 3'b111; end
            18'b110000010100100101: begin rgb_reg = 3'b111; end
            18'b110000010100100110: begin rgb_reg = 3'b111; end
            18'b110000010100100111: begin rgb_reg = 3'b111; end
            18'b110000010100101100: begin rgb_reg = 3'b111; end
            18'b110000010100101101: begin rgb_reg = 3'b111; end
            18'b110000010100111100: begin rgb_reg = 3'b111; end
            18'b110000010100111101: begin rgb_reg = 3'b111; end
            18'b110000011010111110: begin rgb_reg = 3'b111; end
            18'b110000011010111111: begin rgb_reg = 3'b111; end
            18'b110000011011000111: begin rgb_reg = 3'b111; end
            18'b110000011011001000: begin rgb_reg = 3'b111; end
            18'b110000011011001011: begin rgb_reg = 3'b111; end
            18'b110000011011001100: begin rgb_reg = 3'b111; end
            18'b110000011011001101: begin rgb_reg = 3'b111; end
            18'b110000011011010100: begin rgb_reg = 3'b111; end
            18'b110000011011010101: begin rgb_reg = 3'b111; end
            18'b110000011011010110: begin rgb_reg = 3'b111; end
            18'b110000011011011001: begin rgb_reg = 3'b111; end
            18'b110000011011011010: begin rgb_reg = 3'b111; end
            18'b110000011011100010: begin rgb_reg = 3'b111; end
            18'b110000011011100011: begin rgb_reg = 3'b111; end
            18'b110000011011100110: begin rgb_reg = 3'b111; end
            18'b110000011011100111: begin rgb_reg = 3'b111; end
            18'b110000011011101000: begin rgb_reg = 3'b111; end
            18'b110000011011101111: begin rgb_reg = 3'b111; end
            18'b110000011011110000: begin rgb_reg = 3'b111; end
            18'b110000011011110001: begin rgb_reg = 3'b111; end
            18'b110000011011110100: begin rgb_reg = 3'b111; end
            18'b110000011011110101: begin rgb_reg = 3'b111; end
            18'b110000011011111101: begin rgb_reg = 3'b111; end
            18'b110000011011111110: begin rgb_reg = 3'b111; end
            18'b110000011100000001: begin rgb_reg = 3'b111; end
            18'b110000011100000010: begin rgb_reg = 3'b111; end
            18'b110000011100000011: begin rgb_reg = 3'b111; end
            18'b110000011100001111: begin rgb_reg = 3'b111; end
            18'b110000011100010000: begin rgb_reg = 3'b111; end
            18'b110000011100011000: begin rgb_reg = 3'b111; end
            18'b110000011100011001: begin rgb_reg = 3'b111; end
            18'b110000011100100101: begin rgb_reg = 3'b111; end
            18'b110000011100100110: begin rgb_reg = 3'b111; end
            18'b110000011100100111: begin rgb_reg = 3'b111; end
            18'b110000011100101010: begin rgb_reg = 3'b111; end
            18'b110000011100101011: begin rgb_reg = 3'b111; end
            18'b110000011100111100: begin rgb_reg = 3'b111; end
            18'b110000011100111101: begin rgb_reg = 3'b111; end
            18'b110000100010111110: begin rgb_reg = 3'b111; end
            18'b110000100010111111: begin rgb_reg = 3'b111; end
            18'b110000100011000111: begin rgb_reg = 3'b111; end
            18'b110000100011001000: begin rgb_reg = 3'b111; end
            18'b110000100011001011: begin rgb_reg = 3'b111; end
            18'b110000100011001100: begin rgb_reg = 3'b111; end
            18'b110000100011001101: begin rgb_reg = 3'b111; end
            18'b110000100011010100: begin rgb_reg = 3'b111; end
            18'b110000100011010101: begin rgb_reg = 3'b111; end
            18'b110000100011010110: begin rgb_reg = 3'b111; end
            18'b110000100011011001: begin rgb_reg = 3'b111; end
            18'b110000100011011010: begin rgb_reg = 3'b111; end
            18'b110000100011100010: begin rgb_reg = 3'b111; end
            18'b110000100011100011: begin rgb_reg = 3'b111; end
            18'b110000100011100110: begin rgb_reg = 3'b111; end
            18'b110000100011100111: begin rgb_reg = 3'b111; end
            18'b110000100011101000: begin rgb_reg = 3'b111; end
            18'b110000100011101111: begin rgb_reg = 3'b111; end
            18'b110000100011110000: begin rgb_reg = 3'b111; end
            18'b110000100011110001: begin rgb_reg = 3'b111; end
            18'b110000100011110100: begin rgb_reg = 3'b111; end
            18'b110000100011110101: begin rgb_reg = 3'b111; end
            18'b110000100011111101: begin rgb_reg = 3'b111; end
            18'b110000100011111110: begin rgb_reg = 3'b111; end
            18'b110000100100000001: begin rgb_reg = 3'b111; end
            18'b110000100100000010: begin rgb_reg = 3'b111; end
            18'b110000100100000011: begin rgb_reg = 3'b111; end
            18'b110000100100001111: begin rgb_reg = 3'b111; end
            18'b110000100100010000: begin rgb_reg = 3'b111; end
            18'b110000100100011000: begin rgb_reg = 3'b111; end
            18'b110000100100011001: begin rgb_reg = 3'b111; end
            18'b110000100100100101: begin rgb_reg = 3'b111; end
            18'b110000100100100110: begin rgb_reg = 3'b111; end
            18'b110000100100100111: begin rgb_reg = 3'b111; end
            18'b110000100100101010: begin rgb_reg = 3'b111; end
            18'b110000100100101011: begin rgb_reg = 3'b111; end
            18'b110000100100111100: begin rgb_reg = 3'b111; end
            18'b110000100100111101: begin rgb_reg = 3'b111; end
            18'b110000101010111110: begin rgb_reg = 3'b111; end
            18'b110000101010111111: begin rgb_reg = 3'b111; end
            18'b110000101011000000: begin rgb_reg = 3'b111; end
            18'b110000101011000001: begin rgb_reg = 3'b111; end
            18'b110000101011000010: begin rgb_reg = 3'b111; end
            18'b110000101011000011: begin rgb_reg = 3'b111; end
            18'b110000101011000100: begin rgb_reg = 3'b111; end
            18'b110000101011000101: begin rgb_reg = 3'b111; end
            18'b110000101011000110: begin rgb_reg = 3'b111; end
            18'b110000101011000111: begin rgb_reg = 3'b111; end
            18'b110000101011001000: begin rgb_reg = 3'b111; end
            18'b110000101011001100: begin rgb_reg = 3'b111; end
            18'b110000101011001101: begin rgb_reg = 3'b111; end
            18'b110000101011001110: begin rgb_reg = 3'b111; end
            18'b110000101011001111: begin rgb_reg = 3'b111; end
            18'b110000101011010000: begin rgb_reg = 3'b111; end
            18'b110000101011010001: begin rgb_reg = 3'b111; end
            18'b110000101011010010: begin rgb_reg = 3'b111; end
            18'b110000101011010011: begin rgb_reg = 3'b111; end
            18'b110000101011010100: begin rgb_reg = 3'b111; end
            18'b110000101011010101: begin rgb_reg = 3'b111; end
            18'b110000101011011001: begin rgb_reg = 3'b111; end
            18'b110000101011011010: begin rgb_reg = 3'b111; end
            18'b110000101011011011: begin rgb_reg = 3'b111; end
            18'b110000101011011100: begin rgb_reg = 3'b111; end
            18'b110000101011011101: begin rgb_reg = 3'b111; end
            18'b110000101011011110: begin rgb_reg = 3'b111; end
            18'b110000101011011111: begin rgb_reg = 3'b111; end
            18'b110000101011100000: begin rgb_reg = 3'b111; end
            18'b110000101011100001: begin rgb_reg = 3'b111; end
            18'b110000101011100010: begin rgb_reg = 3'b111; end
            18'b110000101011100011: begin rgb_reg = 3'b111; end
            18'b110000101011100111: begin rgb_reg = 3'b111; end
            18'b110000101011101000: begin rgb_reg = 3'b111; end
            18'b110000101011101001: begin rgb_reg = 3'b111; end
            18'b110000101011101010: begin rgb_reg = 3'b111; end
            18'b110000101011101011: begin rgb_reg = 3'b111; end
            18'b110000101011101100: begin rgb_reg = 3'b111; end
            18'b110000101011101101: begin rgb_reg = 3'b111; end
            18'b110000101011101110: begin rgb_reg = 3'b111; end
            18'b110000101011101111: begin rgb_reg = 3'b111; end
            18'b110000101011110000: begin rgb_reg = 3'b111; end
            18'b110000101011110100: begin rgb_reg = 3'b111; end
            18'b110000101011110101: begin rgb_reg = 3'b111; end
            18'b110000101011110110: begin rgb_reg = 3'b111; end
            18'b110000101011110111: begin rgb_reg = 3'b111; end
            18'b110000101011111000: begin rgb_reg = 3'b111; end
            18'b110000101011111001: begin rgb_reg = 3'b111; end
            18'b110000101011111010: begin rgb_reg = 3'b111; end
            18'b110000101011111011: begin rgb_reg = 3'b111; end
            18'b110000101011111100: begin rgb_reg = 3'b111; end
            18'b110000101011111101: begin rgb_reg = 3'b111; end
            18'b110000101011111110: begin rgb_reg = 3'b111; end
            18'b110000101100000001: begin rgb_reg = 3'b111; end
            18'b110000101100000010: begin rgb_reg = 3'b111; end
            18'b110000101100000011: begin rgb_reg = 3'b111; end
            18'b110000101100000100: begin rgb_reg = 3'b111; end
            18'b110000101100000101: begin rgb_reg = 3'b111; end
            18'b110000101100000110: begin rgb_reg = 3'b111; end
            18'b110000101100000111: begin rgb_reg = 3'b111; end
            18'b110000101100001000: begin rgb_reg = 3'b111; end
            18'b110000101100001001: begin rgb_reg = 3'b111; end
            18'b110000101100001010: begin rgb_reg = 3'b111; end
            18'b110000101100001011: begin rgb_reg = 3'b111; end
            18'b110000101100001111: begin rgb_reg = 3'b111; end
            18'b110000101100010000: begin rgb_reg = 3'b111; end
            18'b110000101100010001: begin rgb_reg = 3'b111; end
            18'b110000101100010010: begin rgb_reg = 3'b111; end
            18'b110000101100010011: begin rgb_reg = 3'b111; end
            18'b110000101100010100: begin rgb_reg = 3'b111; end
            18'b110000101100010101: begin rgb_reg = 3'b111; end
            18'b110000101100010110: begin rgb_reg = 3'b111; end
            18'b110000101100010111: begin rgb_reg = 3'b111; end
            18'b110000101100011000: begin rgb_reg = 3'b111; end
            18'b110000101100011001: begin rgb_reg = 3'b111; end
            18'b110000101100100101: begin rgb_reg = 3'b111; end
            18'b110000101100100110: begin rgb_reg = 3'b111; end
            18'b110000101100100111: begin rgb_reg = 3'b111; end
            18'b110000101100101010: begin rgb_reg = 3'b111; end
            18'b110000101100101011: begin rgb_reg = 3'b111; end
            18'b110000101100101100: begin rgb_reg = 3'b111; end
            18'b110000101100101101: begin rgb_reg = 3'b111; end
            18'b110000101100101110: begin rgb_reg = 3'b111; end
            18'b110000101100101111: begin rgb_reg = 3'b111; end
            18'b110000101100110000: begin rgb_reg = 3'b111; end
            18'b110000101100110001: begin rgb_reg = 3'b111; end
            18'b110000101100110010: begin rgb_reg = 3'b111; end
            18'b110000101100110011: begin rgb_reg = 3'b111; end
            18'b110000101100110100: begin rgb_reg = 3'b111; end
            18'b110000101100111000: begin rgb_reg = 3'b111; end
            18'b110000101100111001: begin rgb_reg = 3'b111; end
            18'b110000101100111010: begin rgb_reg = 3'b111; end
            18'b110000101100111011: begin rgb_reg = 3'b111; end
            18'b110000101100111100: begin rgb_reg = 3'b111; end
            18'b110000101100111101: begin rgb_reg = 3'b111; end
            18'b110000101100111110: begin rgb_reg = 3'b111; end
            18'b110000101100111111: begin rgb_reg = 3'b111; end
            18'b110000101101000000: begin rgb_reg = 3'b111; end
            18'b110000101101000001: begin rgb_reg = 3'b111; end
            18'b110000110011000000: begin rgb_reg = 3'b111; end
            18'b110000110011000001: begin rgb_reg = 3'b111; end
            18'b110000110011000010: begin rgb_reg = 3'b111; end
            18'b110000110011000011: begin rgb_reg = 3'b111; end
            18'b110000110011000100: begin rgb_reg = 3'b111; end
            18'b110000110011000101: begin rgb_reg = 3'b111; end
            18'b110000110011000110: begin rgb_reg = 3'b111; end
            18'b110000110011001101: begin rgb_reg = 3'b111; end
            18'b110000110011001110: begin rgb_reg = 3'b111; end
            18'b110000110011001111: begin rgb_reg = 3'b111; end
            18'b110000110011010000: begin rgb_reg = 3'b111; end
            18'b110000110011010001: begin rgb_reg = 3'b111; end
            18'b110000110011010010: begin rgb_reg = 3'b111; end
            18'b110000110011010011: begin rgb_reg = 3'b111; end
            18'b110000110011011011: begin rgb_reg = 3'b111; end
            18'b110000110011011100: begin rgb_reg = 3'b111; end
            18'b110000110011011101: begin rgb_reg = 3'b111; end
            18'b110000110011011110: begin rgb_reg = 3'b111; end
            18'b110000110011011111: begin rgb_reg = 3'b111; end
            18'b110000110011100000: begin rgb_reg = 3'b111; end
            18'b110000110011100001: begin rgb_reg = 3'b111; end
            18'b110000110011101000: begin rgb_reg = 3'b111; end
            18'b110000110011101001: begin rgb_reg = 3'b111; end
            18'b110000110011101010: begin rgb_reg = 3'b111; end
            18'b110000110011101011: begin rgb_reg = 3'b111; end
            18'b110000110011101100: begin rgb_reg = 3'b111; end
            18'b110000110011101101: begin rgb_reg = 3'b111; end
            18'b110000110011101110: begin rgb_reg = 3'b111; end
            18'b110000110011110110: begin rgb_reg = 3'b111; end
            18'b110000110011110111: begin rgb_reg = 3'b111; end
            18'b110000110011111000: begin rgb_reg = 3'b111; end
            18'b110000110011111001: begin rgb_reg = 3'b111; end
            18'b110000110011111010: begin rgb_reg = 3'b111; end
            18'b110000110011111011: begin rgb_reg = 3'b111; end
            18'b110000110011111100: begin rgb_reg = 3'b111; end
            18'b110000110100000001: begin rgb_reg = 3'b111; end
            18'b110000110100000010: begin rgb_reg = 3'b111; end
            18'b110000110100000011: begin rgb_reg = 3'b111; end
            18'b110000110100000100: begin rgb_reg = 3'b111; end
            18'b110000110100000101: begin rgb_reg = 3'b111; end
            18'b110000110100000110: begin rgb_reg = 3'b111; end
            18'b110000110100000111: begin rgb_reg = 3'b111; end
            18'b110000110100001000: begin rgb_reg = 3'b111; end
            18'b110000110100001001: begin rgb_reg = 3'b111; end
            18'b110000110100001010: begin rgb_reg = 3'b111; end
            18'b110000110100001011: begin rgb_reg = 3'b111; end
            18'b110000110100001100: begin rgb_reg = 3'b111; end
            18'b110000110100010001: begin rgb_reg = 3'b111; end
            18'b110000110100010010: begin rgb_reg = 3'b111; end
            18'b110000110100010011: begin rgb_reg = 3'b111; end
            18'b110000110100010100: begin rgb_reg = 3'b111; end
            18'b110000110100010101: begin rgb_reg = 3'b111; end
            18'b110000110100010110: begin rgb_reg = 3'b111; end
            18'b110000110100010111: begin rgb_reg = 3'b111; end
            18'b110000110100100101: begin rgb_reg = 3'b111; end
            18'b110000110100100110: begin rgb_reg = 3'b111; end
            18'b110000110100100111: begin rgb_reg = 3'b111; end
            18'b110000110100101010: begin rgb_reg = 3'b111; end
            18'b110000110100101011: begin rgb_reg = 3'b111; end
            18'b110000110100101100: begin rgb_reg = 3'b111; end
            18'b110000110100101101: begin rgb_reg = 3'b111; end
            18'b110000110100101110: begin rgb_reg = 3'b111; end
            18'b110000110100101111: begin rgb_reg = 3'b111; end
            18'b110000110100110000: begin rgb_reg = 3'b111; end
            18'b110000110100110001: begin rgb_reg = 3'b111; end
            18'b110000110100110010: begin rgb_reg = 3'b111; end
            18'b110000110100110011: begin rgb_reg = 3'b111; end
            18'b110000110100110100: begin rgb_reg = 3'b111; end
            18'b110000110100110111: begin rgb_reg = 3'b111; end
            18'b110000110100111000: begin rgb_reg = 3'b111; end
            18'b110000110100111001: begin rgb_reg = 3'b111; end
            18'b110000110100111010: begin rgb_reg = 3'b111; end
            18'b110000110100111011: begin rgb_reg = 3'b111; end
            18'b110000110100111100: begin rgb_reg = 3'b111; end
            18'b110000110100111101: begin rgb_reg = 3'b111; end
            18'b110000110100111110: begin rgb_reg = 3'b111; end
            18'b110000110100111111: begin rgb_reg = 3'b111; end
            18'b110000110101000000: begin rgb_reg = 3'b111; end
            18'b110000110101000001: begin rgb_reg = 3'b111; end
            18'b110000110101000010: begin rgb_reg = 3'b111; end
            18'b110000111011000000: begin rgb_reg = 3'b111; end
            18'b110000111011000001: begin rgb_reg = 3'b111; end
            18'b110000111011000010: begin rgb_reg = 3'b111; end
            18'b110000111011000011: begin rgb_reg = 3'b111; end
            18'b110000111011000100: begin rgb_reg = 3'b111; end
            18'b110000111011000101: begin rgb_reg = 3'b111; end
            18'b110000111011000110: begin rgb_reg = 3'b111; end
            18'b110000111011001110: begin rgb_reg = 3'b111; end
            18'b110000111011001111: begin rgb_reg = 3'b111; end
            18'b110000111011010000: begin rgb_reg = 3'b111; end
            18'b110000111011010001: begin rgb_reg = 3'b111; end
            18'b110000111011010010: begin rgb_reg = 3'b111; end
            18'b110000111011010011: begin rgb_reg = 3'b111; end
            18'b110000111011011011: begin rgb_reg = 3'b111; end
            18'b110000111011011100: begin rgb_reg = 3'b111; end
            18'b110000111011011101: begin rgb_reg = 3'b111; end
            18'b110000111011011110: begin rgb_reg = 3'b111; end
            18'b110000111011011111: begin rgb_reg = 3'b111; end
            18'b110000111011100000: begin rgb_reg = 3'b111; end
            18'b110000111011100001: begin rgb_reg = 3'b111; end
            18'b110000111011101001: begin rgb_reg = 3'b111; end
            18'b110000111011101010: begin rgb_reg = 3'b111; end
            18'b110000111011101011: begin rgb_reg = 3'b111; end
            18'b110000111011101100: begin rgb_reg = 3'b111; end
            18'b110000111011101101: begin rgb_reg = 3'b111; end
            18'b110000111011101110: begin rgb_reg = 3'b111; end
            18'b110000111011110110: begin rgb_reg = 3'b111; end
            18'b110000111011110111: begin rgb_reg = 3'b111; end
            18'b110000111011111000: begin rgb_reg = 3'b111; end
            18'b110000111011111001: begin rgb_reg = 3'b111; end
            18'b110000111011111010: begin rgb_reg = 3'b111; end
            18'b110000111011111011: begin rgb_reg = 3'b111; end
            18'b110000111011111100: begin rgb_reg = 3'b111; end
            18'b110000111100000001: begin rgb_reg = 3'b111; end
            18'b110000111100000010: begin rgb_reg = 3'b111; end
            18'b110000111100000011: begin rgb_reg = 3'b111; end
            18'b110000111100000100: begin rgb_reg = 3'b111; end
            18'b110000111100000101: begin rgb_reg = 3'b111; end
            18'b110000111100000110: begin rgb_reg = 3'b111; end
            18'b110000111100000111: begin rgb_reg = 3'b111; end
            18'b110000111100001000: begin rgb_reg = 3'b111; end
            18'b110000111100001001: begin rgb_reg = 3'b111; end
            18'b110000111100001010: begin rgb_reg = 3'b111; end
            18'b110000111100001011: begin rgb_reg = 3'b111; end
            18'b110000111100010001: begin rgb_reg = 3'b111; end
            18'b110000111100010010: begin rgb_reg = 3'b111; end
            18'b110000111100010011: begin rgb_reg = 3'b111; end
            18'b110000111100010100: begin rgb_reg = 3'b111; end
            18'b110000111100010101: begin rgb_reg = 3'b111; end
            18'b110000111100010110: begin rgb_reg = 3'b111; end
            18'b110000111100010111: begin rgb_reg = 3'b111; end
            18'b110000111100100101: begin rgb_reg = 3'b111; end
            18'b110000111100100110: begin rgb_reg = 3'b111; end
            18'b110000111100101010: begin rgb_reg = 3'b111; end
            18'b110000111100101011: begin rgb_reg = 3'b111; end
            18'b110000111100101100: begin rgb_reg = 3'b111; end
            18'b110000111100101101: begin rgb_reg = 3'b111; end
            18'b110000111100101110: begin rgb_reg = 3'b111; end
            18'b110000111100101111: begin rgb_reg = 3'b111; end
            18'b110000111100110000: begin rgb_reg = 3'b111; end
            18'b110000111100110001: begin rgb_reg = 3'b111; end
            18'b110000111100110010: begin rgb_reg = 3'b111; end
            18'b110000111100110011: begin rgb_reg = 3'b111; end
            18'b110000111100110100: begin rgb_reg = 3'b111; end
            18'b110000111100110111: begin rgb_reg = 3'b111; end
            18'b110000111100111000: begin rgb_reg = 3'b111; end
            18'b110000111100111001: begin rgb_reg = 3'b111; end
            18'b110000111100111010: begin rgb_reg = 3'b111; end
            18'b110000111100111011: begin rgb_reg = 3'b111; end
            18'b110000111100111100: begin rgb_reg = 3'b111; end
            18'b110000111100111101: begin rgb_reg = 3'b111; end
            18'b110000111100111110: begin rgb_reg = 3'b111; end
            18'b110000111100111111: begin rgb_reg = 3'b111; end
            18'b110000111101000000: begin rgb_reg = 3'b111; end
            18'b110000111101000001: begin rgb_reg = 3'b111; end
            18'b110001110010011000: begin rgb_reg = 3'b111; end
            18'b110001110010011001: begin rgb_reg = 3'b111; end
            18'b110001110010100000: begin rgb_reg = 3'b111; end
            18'b110001110010100001: begin rgb_reg = 3'b111; end
            18'b110001110010111100: begin rgb_reg = 3'b111; end
            18'b110001110010111101: begin rgb_reg = 3'b111; end
            18'b110001110011011000: begin rgb_reg = 3'b111; end
            18'b110001110011011001: begin rgb_reg = 3'b111; end
            18'b110001110011011010: begin rgb_reg = 3'b111; end
            18'b110001110011011011: begin rgb_reg = 3'b111; end
            18'b110001110011011100: begin rgb_reg = 3'b111; end
            18'b110001110011011101: begin rgb_reg = 3'b111; end
            18'b110001110011011110: begin rgb_reg = 3'b111; end
            18'b110001110011011111: begin rgb_reg = 3'b111; end
            18'b110001110011100000: begin rgb_reg = 3'b111; end
            18'b110001110011100001: begin rgb_reg = 3'b111; end
            18'b110001110011111100: begin rgb_reg = 3'b111; end
            18'b110001110011111101: begin rgb_reg = 3'b111; end
            18'b110001110101001110: begin rgb_reg = 3'b111; end
            18'b110001110101001111: begin rgb_reg = 3'b111; end
            18'b110001110101011110: begin rgb_reg = 3'b111; end
            18'b110001110101011111: begin rgb_reg = 3'b111; end
            18'b110001111010011000: begin rgb_reg = 3'b111; end
            18'b110001111010011001: begin rgb_reg = 3'b111; end
            18'b110001111010100000: begin rgb_reg = 3'b111; end
            18'b110001111010100001: begin rgb_reg = 3'b111; end
            18'b110001111010111100: begin rgb_reg = 3'b111; end
            18'b110001111010111101: begin rgb_reg = 3'b111; end
            18'b110001111011011000: begin rgb_reg = 3'b111; end
            18'b110001111011011001: begin rgb_reg = 3'b111; end
            18'b110001111011011010: begin rgb_reg = 3'b111; end
            18'b110001111011011011: begin rgb_reg = 3'b111; end
            18'b110001111011011100: begin rgb_reg = 3'b111; end
            18'b110001111011011101: begin rgb_reg = 3'b111; end
            18'b110001111011011110: begin rgb_reg = 3'b111; end
            18'b110001111011011111: begin rgb_reg = 3'b111; end
            18'b110001111011100000: begin rgb_reg = 3'b111; end
            18'b110001111011100001: begin rgb_reg = 3'b111; end
            18'b110001111011111100: begin rgb_reg = 3'b111; end
            18'b110001111011111101: begin rgb_reg = 3'b111; end
            18'b110001111101001110: begin rgb_reg = 3'b111; end
            18'b110001111101001111: begin rgb_reg = 3'b111; end
            18'b110001111101011110: begin rgb_reg = 3'b111; end
            18'b110001111101011111: begin rgb_reg = 3'b111; end
            18'b110010000010011000: begin rgb_reg = 3'b111; end
            18'b110010000010011001: begin rgb_reg = 3'b111; end
            18'b110010000010011010: begin rgb_reg = 3'b111; end
            18'b110010000010011011: begin rgb_reg = 3'b111; end
            18'b110010000010100000: begin rgb_reg = 3'b111; end
            18'b110010000010100001: begin rgb_reg = 3'b111; end
            18'b110010000011011100: begin rgb_reg = 3'b111; end
            18'b110010000011011101: begin rgb_reg = 3'b111; end
            18'b110010000011111100: begin rgb_reg = 3'b111; end
            18'b110010000011111101: begin rgb_reg = 3'b111; end
            18'b110010000101011110: begin rgb_reg = 3'b111; end
            18'b110010000101011111: begin rgb_reg = 3'b111; end
            18'b110010001010011000: begin rgb_reg = 3'b111; end
            18'b110010001010011001: begin rgb_reg = 3'b111; end
            18'b110010001010011010: begin rgb_reg = 3'b111; end
            18'b110010001010011011: begin rgb_reg = 3'b111; end
            18'b110010001010100000: begin rgb_reg = 3'b111; end
            18'b110010001010100001: begin rgb_reg = 3'b111; end
            18'b110010001011011100: begin rgb_reg = 3'b111; end
            18'b110010001011011101: begin rgb_reg = 3'b111; end
            18'b110010001011111100: begin rgb_reg = 3'b111; end
            18'b110010001011111101: begin rgb_reg = 3'b111; end
            18'b110010001101011110: begin rgb_reg = 3'b111; end
            18'b110010001101011111: begin rgb_reg = 3'b111; end
            18'b110010010010011000: begin rgb_reg = 3'b111; end
            18'b110010010010011001: begin rgb_reg = 3'b111; end
            18'b110010010010011100: begin rgb_reg = 3'b111; end
            18'b110010010010011101: begin rgb_reg = 3'b111; end
            18'b110010010010100000: begin rgb_reg = 3'b111; end
            18'b110010010010100001: begin rgb_reg = 3'b111; end
            18'b110010010010100110: begin rgb_reg = 3'b111; end
            18'b110010010010100111: begin rgb_reg = 3'b111; end
            18'b110010010010101000: begin rgb_reg = 3'b111; end
            18'b110010010010101001: begin rgb_reg = 3'b111; end
            18'b110010010010101010: begin rgb_reg = 3'b111; end
            18'b110010010010101011: begin rgb_reg = 3'b111; end
            18'b110010010010110000: begin rgb_reg = 3'b111; end
            18'b110010010010110001: begin rgb_reg = 3'b111; end
            18'b110010010010110100: begin rgb_reg = 3'b111; end
            18'b110010010010110101: begin rgb_reg = 3'b111; end
            18'b110010010010110110: begin rgb_reg = 3'b111; end
            18'b110010010010110111: begin rgb_reg = 3'b111; end
            18'b110010010010111100: begin rgb_reg = 3'b111; end
            18'b110010010010111101: begin rgb_reg = 3'b111; end
            18'b110010010011000000: begin rgb_reg = 3'b111; end
            18'b110010010011000001: begin rgb_reg = 3'b111; end
            18'b110010010011000010: begin rgb_reg = 3'b111; end
            18'b110010010011000011: begin rgb_reg = 3'b111; end
            18'b110010010011000100: begin rgb_reg = 3'b111; end
            18'b110010010011000101: begin rgb_reg = 3'b111; end
            18'b110010010011000110: begin rgb_reg = 3'b111; end
            18'b110010010011000111: begin rgb_reg = 3'b111; end
            18'b110010010011011100: begin rgb_reg = 3'b111; end
            18'b110010010011011101: begin rgb_reg = 3'b111; end
            18'b110010010011100100: begin rgb_reg = 3'b111; end
            18'b110010010011100101: begin rgb_reg = 3'b111; end
            18'b110010010011101000: begin rgb_reg = 3'b111; end
            18'b110010010011101001: begin rgb_reg = 3'b111; end
            18'b110010010011101010: begin rgb_reg = 3'b111; end
            18'b110010010011101011: begin rgb_reg = 3'b111; end
            18'b110010010011110010: begin rgb_reg = 3'b111; end
            18'b110010010011110011: begin rgb_reg = 3'b111; end
            18'b110010010011110100: begin rgb_reg = 3'b111; end
            18'b110010010011110101: begin rgb_reg = 3'b111; end
            18'b110010010011110110: begin rgb_reg = 3'b111; end
            18'b110010010011110111: begin rgb_reg = 3'b111; end
            18'b110010010011111100: begin rgb_reg = 3'b111; end
            18'b110010010011111101: begin rgb_reg = 3'b111; end
            18'b110010010100000010: begin rgb_reg = 3'b111; end
            18'b110010010100000011: begin rgb_reg = 3'b111; end
            18'b110010010100001000: begin rgb_reg = 3'b111; end
            18'b110010010100001001: begin rgb_reg = 3'b111; end
            18'b110010010100001010: begin rgb_reg = 3'b111; end
            18'b110010010100001011: begin rgb_reg = 3'b111; end
            18'b110010010100001100: begin rgb_reg = 3'b111; end
            18'b110010010100001101: begin rgb_reg = 3'b111; end
            18'b110010010100010010: begin rgb_reg = 3'b111; end
            18'b110010010100010011: begin rgb_reg = 3'b111; end
            18'b110010010100010110: begin rgb_reg = 3'b111; end
            18'b110010010100010111: begin rgb_reg = 3'b111; end
            18'b110010010100011000: begin rgb_reg = 3'b111; end
            18'b110010010100011001: begin rgb_reg = 3'b111; end
            18'b110010010100011110: begin rgb_reg = 3'b111; end
            18'b110010010100011111: begin rgb_reg = 3'b111; end
            18'b110010010100100000: begin rgb_reg = 3'b111; end
            18'b110010010100100001: begin rgb_reg = 3'b111; end
            18'b110010010100100010: begin rgb_reg = 3'b111; end
            18'b110010010100100011: begin rgb_reg = 3'b111; end
            18'b110010010100100100: begin rgb_reg = 3'b111; end
            18'b110010010100100101: begin rgb_reg = 3'b111; end
            18'b110010010100101010: begin rgb_reg = 3'b111; end
            18'b110010010100101011: begin rgb_reg = 3'b111; end
            18'b110010010100110010: begin rgb_reg = 3'b111; end
            18'b110010010100110011: begin rgb_reg = 3'b111; end
            18'b110010010100111000: begin rgb_reg = 3'b111; end
            18'b110010010100111001: begin rgb_reg = 3'b111; end
            18'b110010010100111010: begin rgb_reg = 3'b111; end
            18'b110010010100111011: begin rgb_reg = 3'b111; end
            18'b110010010100111100: begin rgb_reg = 3'b111; end
            18'b110010010100111101: begin rgb_reg = 3'b111; end
            18'b110010010101000010: begin rgb_reg = 3'b111; end
            18'b110010010101000011: begin rgb_reg = 3'b111; end
            18'b110010010101000100: begin rgb_reg = 3'b111; end
            18'b110010010101000101: begin rgb_reg = 3'b111; end
            18'b110010010101000110: begin rgb_reg = 3'b111; end
            18'b110010010101000111: begin rgb_reg = 3'b111; end
            18'b110010010101001000: begin rgb_reg = 3'b111; end
            18'b110010010101001001: begin rgb_reg = 3'b111; end
            18'b110010010101001110: begin rgb_reg = 3'b111; end
            18'b110010010101001111: begin rgb_reg = 3'b111; end
            18'b110010010101010100: begin rgb_reg = 3'b111; end
            18'b110010010101010101: begin rgb_reg = 3'b111; end
            18'b110010010101010110: begin rgb_reg = 3'b111; end
            18'b110010010101010111: begin rgb_reg = 3'b111; end
            18'b110010010101011000: begin rgb_reg = 3'b111; end
            18'b110010010101011001: begin rgb_reg = 3'b111; end
            18'b110010010101011110: begin rgb_reg = 3'b111; end
            18'b110010010101011111: begin rgb_reg = 3'b111; end
            18'b110010010101100010: begin rgb_reg = 3'b111; end
            18'b110010010101100011: begin rgb_reg = 3'b111; end
            18'b110010010101100100: begin rgb_reg = 3'b111; end
            18'b110010010101100101: begin rgb_reg = 3'b111; end
            18'b110010011010011000: begin rgb_reg = 3'b111; end
            18'b110010011010011001: begin rgb_reg = 3'b111; end
            18'b110010011010011100: begin rgb_reg = 3'b111; end
            18'b110010011010011101: begin rgb_reg = 3'b111; end
            18'b110010011010100000: begin rgb_reg = 3'b111; end
            18'b110010011010100001: begin rgb_reg = 3'b111; end
            18'b110010011010100110: begin rgb_reg = 3'b111; end
            18'b110010011010100111: begin rgb_reg = 3'b111; end
            18'b110010011010101000: begin rgb_reg = 3'b111; end
            18'b110010011010101001: begin rgb_reg = 3'b111; end
            18'b110010011010101010: begin rgb_reg = 3'b111; end
            18'b110010011010101011: begin rgb_reg = 3'b111; end
            18'b110010011010110000: begin rgb_reg = 3'b111; end
            18'b110010011010110001: begin rgb_reg = 3'b111; end
            18'b110010011010110100: begin rgb_reg = 3'b111; end
            18'b110010011010110101: begin rgb_reg = 3'b111; end
            18'b110010011010110110: begin rgb_reg = 3'b111; end
            18'b110010011010110111: begin rgb_reg = 3'b111; end
            18'b110010011010111100: begin rgb_reg = 3'b111; end
            18'b110010011010111101: begin rgb_reg = 3'b111; end
            18'b110010011011000000: begin rgb_reg = 3'b111; end
            18'b110010011011000001: begin rgb_reg = 3'b111; end
            18'b110010011011000010: begin rgb_reg = 3'b111; end
            18'b110010011011000011: begin rgb_reg = 3'b111; end
            18'b110010011011000100: begin rgb_reg = 3'b111; end
            18'b110010011011000101: begin rgb_reg = 3'b111; end
            18'b110010011011000110: begin rgb_reg = 3'b111; end
            18'b110010011011000111: begin rgb_reg = 3'b111; end
            18'b110010011011011100: begin rgb_reg = 3'b111; end
            18'b110010011011011101: begin rgb_reg = 3'b111; end
            18'b110010011011100100: begin rgb_reg = 3'b111; end
            18'b110010011011100101: begin rgb_reg = 3'b111; end
            18'b110010011011101000: begin rgb_reg = 3'b111; end
            18'b110010011011101001: begin rgb_reg = 3'b111; end
            18'b110010011011101010: begin rgb_reg = 3'b111; end
            18'b110010011011101011: begin rgb_reg = 3'b111; end
            18'b110010011011110010: begin rgb_reg = 3'b111; end
            18'b110010011011110011: begin rgb_reg = 3'b111; end
            18'b110010011011110100: begin rgb_reg = 3'b111; end
            18'b110010011011110101: begin rgb_reg = 3'b111; end
            18'b110010011011110110: begin rgb_reg = 3'b111; end
            18'b110010011011110111: begin rgb_reg = 3'b111; end
            18'b110010011011111100: begin rgb_reg = 3'b111; end
            18'b110010011011111101: begin rgb_reg = 3'b111; end
            18'b110010011100000010: begin rgb_reg = 3'b111; end
            18'b110010011100000011: begin rgb_reg = 3'b111; end
            18'b110010011100001000: begin rgb_reg = 3'b111; end
            18'b110010011100001001: begin rgb_reg = 3'b111; end
            18'b110010011100001010: begin rgb_reg = 3'b111; end
            18'b110010011100001011: begin rgb_reg = 3'b111; end
            18'b110010011100001100: begin rgb_reg = 3'b111; end
            18'b110010011100001101: begin rgb_reg = 3'b111; end
            18'b110010011100010010: begin rgb_reg = 3'b111; end
            18'b110010011100010011: begin rgb_reg = 3'b111; end
            18'b110010011100010110: begin rgb_reg = 3'b111; end
            18'b110010011100010111: begin rgb_reg = 3'b111; end
            18'b110010011100011000: begin rgb_reg = 3'b111; end
            18'b110010011100011001: begin rgb_reg = 3'b111; end
            18'b110010011100011110: begin rgb_reg = 3'b111; end
            18'b110010011100011111: begin rgb_reg = 3'b111; end
            18'b110010011100100000: begin rgb_reg = 3'b111; end
            18'b110010011100100001: begin rgb_reg = 3'b111; end
            18'b110010011100100010: begin rgb_reg = 3'b111; end
            18'b110010011100100011: begin rgb_reg = 3'b111; end
            18'b110010011100100100: begin rgb_reg = 3'b111; end
            18'b110010011100100101: begin rgb_reg = 3'b111; end
            18'b110010011100101010: begin rgb_reg = 3'b111; end
            18'b110010011100101011: begin rgb_reg = 3'b111; end
            18'b110010011100110010: begin rgb_reg = 3'b111; end
            18'b110010011100110011: begin rgb_reg = 3'b111; end
            18'b110010011100111000: begin rgb_reg = 3'b111; end
            18'b110010011100111001: begin rgb_reg = 3'b111; end
            18'b110010011100111010: begin rgb_reg = 3'b111; end
            18'b110010011100111011: begin rgb_reg = 3'b111; end
            18'b110010011100111100: begin rgb_reg = 3'b111; end
            18'b110010011100111101: begin rgb_reg = 3'b111; end
            18'b110010011101000010: begin rgb_reg = 3'b111; end
            18'b110010011101000011: begin rgb_reg = 3'b111; end
            18'b110010011101000100: begin rgb_reg = 3'b111; end
            18'b110010011101000101: begin rgb_reg = 3'b111; end
            18'b110010011101000110: begin rgb_reg = 3'b111; end
            18'b110010011101000111: begin rgb_reg = 3'b111; end
            18'b110010011101001000: begin rgb_reg = 3'b111; end
            18'b110010011101001001: begin rgb_reg = 3'b111; end
            18'b110010011101001110: begin rgb_reg = 3'b111; end
            18'b110010011101001111: begin rgb_reg = 3'b111; end
            18'b110010011101010100: begin rgb_reg = 3'b111; end
            18'b110010011101010101: begin rgb_reg = 3'b111; end
            18'b110010011101010110: begin rgb_reg = 3'b111; end
            18'b110010011101010111: begin rgb_reg = 3'b111; end
            18'b110010011101011000: begin rgb_reg = 3'b111; end
            18'b110010011101011001: begin rgb_reg = 3'b111; end
            18'b110010011101011110: begin rgb_reg = 3'b111; end
            18'b110010011101011111: begin rgb_reg = 3'b111; end
            18'b110010011101100010: begin rgb_reg = 3'b111; end
            18'b110010011101100011: begin rgb_reg = 3'b111; end
            18'b110010011101100100: begin rgb_reg = 3'b111; end
            18'b110010011101100101: begin rgb_reg = 3'b111; end
            18'b110010100010011000: begin rgb_reg = 3'b111; end
            18'b110010100010011001: begin rgb_reg = 3'b111; end
            18'b110010100010011110: begin rgb_reg = 3'b111; end
            18'b110010100010011111: begin rgb_reg = 3'b111; end
            18'b110010100010100000: begin rgb_reg = 3'b111; end
            18'b110010100010100001: begin rgb_reg = 3'b111; end
            18'b110010100010101100: begin rgb_reg = 3'b111; end
            18'b110010100010101101: begin rgb_reg = 3'b111; end
            18'b110010100010110000: begin rgb_reg = 3'b111; end
            18'b110010100010110001: begin rgb_reg = 3'b111; end
            18'b110010100010110010: begin rgb_reg = 3'b111; end
            18'b110010100010110011: begin rgb_reg = 3'b111; end
            18'b110010100010111000: begin rgb_reg = 3'b111; end
            18'b110010100010111001: begin rgb_reg = 3'b111; end
            18'b110010100010111100: begin rgb_reg = 3'b111; end
            18'b110010100010111101: begin rgb_reg = 3'b111; end
            18'b110010100011000000: begin rgb_reg = 3'b111; end
            18'b110010100011000001: begin rgb_reg = 3'b111; end
            18'b110010100011001000: begin rgb_reg = 3'b111; end
            18'b110010100011001001: begin rgb_reg = 3'b111; end
            18'b110010100011011100: begin rgb_reg = 3'b111; end
            18'b110010100011011101: begin rgb_reg = 3'b111; end
            18'b110010100011100100: begin rgb_reg = 3'b111; end
            18'b110010100011100101: begin rgb_reg = 3'b111; end
            18'b110010100011100110: begin rgb_reg = 3'b111; end
            18'b110010100011100111: begin rgb_reg = 3'b111; end
            18'b110010100011101100: begin rgb_reg = 3'b111; end
            18'b110010100011101101: begin rgb_reg = 3'b111; end
            18'b110010100011111000: begin rgb_reg = 3'b111; end
            18'b110010100011111001: begin rgb_reg = 3'b111; end
            18'b110010100011111100: begin rgb_reg = 3'b111; end
            18'b110010100011111101: begin rgb_reg = 3'b111; end
            18'b110010100100000000: begin rgb_reg = 3'b111; end
            18'b110010100100000001: begin rgb_reg = 3'b111; end
            18'b110010100100001110: begin rgb_reg = 3'b111; end
            18'b110010100100001111: begin rgb_reg = 3'b111; end
            18'b110010100100010010: begin rgb_reg = 3'b111; end
            18'b110010100100010011: begin rgb_reg = 3'b111; end
            18'b110010100100010100: begin rgb_reg = 3'b111; end
            18'b110010100100010101: begin rgb_reg = 3'b111; end
            18'b110010100100011010: begin rgb_reg = 3'b111; end
            18'b110010100100011011: begin rgb_reg = 3'b111; end
            18'b110010100100011110: begin rgb_reg = 3'b111; end
            18'b110010100100011111: begin rgb_reg = 3'b111; end
            18'b110010100100100110: begin rgb_reg = 3'b111; end
            18'b110010100100100111: begin rgb_reg = 3'b111; end
            18'b110010100100101010: begin rgb_reg = 3'b111; end
            18'b110010100100101011: begin rgb_reg = 3'b111; end
            18'b110010100100110010: begin rgb_reg = 3'b111; end
            18'b110010100100110011: begin rgb_reg = 3'b111; end
            18'b110010100100111110: begin rgb_reg = 3'b111; end
            18'b110010100100111111: begin rgb_reg = 3'b111; end
            18'b110010100101000010: begin rgb_reg = 3'b111; end
            18'b110010100101000011: begin rgb_reg = 3'b111; end
            18'b110010100101001010: begin rgb_reg = 3'b111; end
            18'b110010100101001011: begin rgb_reg = 3'b111; end
            18'b110010100101001110: begin rgb_reg = 3'b111; end
            18'b110010100101001111: begin rgb_reg = 3'b111; end
            18'b110010100101010010: begin rgb_reg = 3'b111; end
            18'b110010100101010011: begin rgb_reg = 3'b111; end
            18'b110010100101011010: begin rgb_reg = 3'b111; end
            18'b110010100101011011: begin rgb_reg = 3'b111; end
            18'b110010100101011110: begin rgb_reg = 3'b111; end
            18'b110010100101011111: begin rgb_reg = 3'b111; end
            18'b110010100101100000: begin rgb_reg = 3'b111; end
            18'b110010100101100001: begin rgb_reg = 3'b111; end
            18'b110010100101100110: begin rgb_reg = 3'b111; end
            18'b110010100101100111: begin rgb_reg = 3'b111; end
            18'b110010101010011000: begin rgb_reg = 3'b111; end
            18'b110010101010011001: begin rgb_reg = 3'b111; end
            18'b110010101010011110: begin rgb_reg = 3'b111; end
            18'b110010101010011111: begin rgb_reg = 3'b111; end
            18'b110010101010100000: begin rgb_reg = 3'b111; end
            18'b110010101010100001: begin rgb_reg = 3'b111; end
            18'b110010101010101100: begin rgb_reg = 3'b111; end
            18'b110010101010101101: begin rgb_reg = 3'b111; end
            18'b110010101010110000: begin rgb_reg = 3'b111; end
            18'b110010101010110001: begin rgb_reg = 3'b111; end
            18'b110010101010110010: begin rgb_reg = 3'b111; end
            18'b110010101010110011: begin rgb_reg = 3'b111; end
            18'b110010101010111000: begin rgb_reg = 3'b111; end
            18'b110010101010111001: begin rgb_reg = 3'b111; end
            18'b110010101010111100: begin rgb_reg = 3'b111; end
            18'b110010101010111101: begin rgb_reg = 3'b111; end
            18'b110010101011000000: begin rgb_reg = 3'b111; end
            18'b110010101011000001: begin rgb_reg = 3'b111; end
            18'b110010101011001000: begin rgb_reg = 3'b111; end
            18'b110010101011001001: begin rgb_reg = 3'b111; end
            18'b110010101011011100: begin rgb_reg = 3'b111; end
            18'b110010101011011101: begin rgb_reg = 3'b111; end
            18'b110010101011100100: begin rgb_reg = 3'b111; end
            18'b110010101011100101: begin rgb_reg = 3'b111; end
            18'b110010101011100110: begin rgb_reg = 3'b111; end
            18'b110010101011100111: begin rgb_reg = 3'b111; end
            18'b110010101011101100: begin rgb_reg = 3'b111; end
            18'b110010101011101101: begin rgb_reg = 3'b111; end
            18'b110010101011111000: begin rgb_reg = 3'b111; end
            18'b110010101011111001: begin rgb_reg = 3'b111; end
            18'b110010101011111100: begin rgb_reg = 3'b111; end
            18'b110010101011111101: begin rgb_reg = 3'b111; end
            18'b110010101100000000: begin rgb_reg = 3'b111; end
            18'b110010101100000001: begin rgb_reg = 3'b111; end
            18'b110010101100001110: begin rgb_reg = 3'b111; end
            18'b110010101100001111: begin rgb_reg = 3'b111; end
            18'b110010101100010010: begin rgb_reg = 3'b111; end
            18'b110010101100010011: begin rgb_reg = 3'b111; end
            18'b110010101100010100: begin rgb_reg = 3'b111; end
            18'b110010101100010101: begin rgb_reg = 3'b111; end
            18'b110010101100011010: begin rgb_reg = 3'b111; end
            18'b110010101100011011: begin rgb_reg = 3'b111; end
            18'b110010101100011110: begin rgb_reg = 3'b111; end
            18'b110010101100011111: begin rgb_reg = 3'b111; end
            18'b110010101100100110: begin rgb_reg = 3'b111; end
            18'b110010101100100111: begin rgb_reg = 3'b111; end
            18'b110010101100101010: begin rgb_reg = 3'b111; end
            18'b110010101100101011: begin rgb_reg = 3'b111; end
            18'b110010101100110010: begin rgb_reg = 3'b111; end
            18'b110010101100110011: begin rgb_reg = 3'b111; end
            18'b110010101100111110: begin rgb_reg = 3'b111; end
            18'b110010101100111111: begin rgb_reg = 3'b111; end
            18'b110010101101000010: begin rgb_reg = 3'b111; end
            18'b110010101101000011: begin rgb_reg = 3'b111; end
            18'b110010101101001010: begin rgb_reg = 3'b111; end
            18'b110010101101001011: begin rgb_reg = 3'b111; end
            18'b110010101101001110: begin rgb_reg = 3'b111; end
            18'b110010101101001111: begin rgb_reg = 3'b111; end
            18'b110010101101010010: begin rgb_reg = 3'b111; end
            18'b110010101101010011: begin rgb_reg = 3'b111; end
            18'b110010101101011010: begin rgb_reg = 3'b111; end
            18'b110010101101011011: begin rgb_reg = 3'b111; end
            18'b110010101101011110: begin rgb_reg = 3'b111; end
            18'b110010101101011111: begin rgb_reg = 3'b111; end
            18'b110010101101100000: begin rgb_reg = 3'b111; end
            18'b110010101101100001: begin rgb_reg = 3'b111; end
            18'b110010101101100110: begin rgb_reg = 3'b111; end
            18'b110010101101100111: begin rgb_reg = 3'b111; end
            18'b110010110010011000: begin rgb_reg = 3'b111; end
            18'b110010110010011001: begin rgb_reg = 3'b111; end
            18'b110010110010100000: begin rgb_reg = 3'b111; end
            18'b110010110010100001: begin rgb_reg = 3'b111; end
            18'b110010110010100110: begin rgb_reg = 3'b111; end
            18'b110010110010100111: begin rgb_reg = 3'b111; end
            18'b110010110010101000: begin rgb_reg = 3'b111; end
            18'b110010110010101001: begin rgb_reg = 3'b111; end
            18'b110010110010101010: begin rgb_reg = 3'b111; end
            18'b110010110010101011: begin rgb_reg = 3'b111; end
            18'b110010110010101100: begin rgb_reg = 3'b111; end
            18'b110010110010101101: begin rgb_reg = 3'b111; end
            18'b110010110010110000: begin rgb_reg = 3'b111; end
            18'b110010110010110001: begin rgb_reg = 3'b111; end
            18'b110010110010111100: begin rgb_reg = 3'b111; end
            18'b110010110010111101: begin rgb_reg = 3'b111; end
            18'b110010110011000000: begin rgb_reg = 3'b111; end
            18'b110010110011000001: begin rgb_reg = 3'b111; end
            18'b110010110011001000: begin rgb_reg = 3'b111; end
            18'b110010110011001001: begin rgb_reg = 3'b111; end
            18'b110010110011011100: begin rgb_reg = 3'b111; end
            18'b110010110011011101: begin rgb_reg = 3'b111; end
            18'b110010110011100100: begin rgb_reg = 3'b111; end
            18'b110010110011100101: begin rgb_reg = 3'b111; end
            18'b110010110011110010: begin rgb_reg = 3'b111; end
            18'b110010110011110011: begin rgb_reg = 3'b111; end
            18'b110010110011110100: begin rgb_reg = 3'b111; end
            18'b110010110011110101: begin rgb_reg = 3'b111; end
            18'b110010110011110110: begin rgb_reg = 3'b111; end
            18'b110010110011110111: begin rgb_reg = 3'b111; end
            18'b110010110011111000: begin rgb_reg = 3'b111; end
            18'b110010110011111001: begin rgb_reg = 3'b111; end
            18'b110010110011111100: begin rgb_reg = 3'b111; end
            18'b110010110011111101: begin rgb_reg = 3'b111; end
            18'b110010110011111110: begin rgb_reg = 3'b111; end
            18'b110010110011111111: begin rgb_reg = 3'b111; end
            18'b110010110100001000: begin rgb_reg = 3'b111; end
            18'b110010110100001001: begin rgb_reg = 3'b111; end
            18'b110010110100001010: begin rgb_reg = 3'b111; end
            18'b110010110100001011: begin rgb_reg = 3'b111; end
            18'b110010110100001100: begin rgb_reg = 3'b111; end
            18'b110010110100001101: begin rgb_reg = 3'b111; end
            18'b110010110100001110: begin rgb_reg = 3'b111; end
            18'b110010110100001111: begin rgb_reg = 3'b111; end
            18'b110010110100010010: begin rgb_reg = 3'b111; end
            18'b110010110100010011: begin rgb_reg = 3'b111; end
            18'b110010110100011110: begin rgb_reg = 3'b111; end
            18'b110010110100011111: begin rgb_reg = 3'b111; end
            18'b110010110100100110: begin rgb_reg = 3'b111; end
            18'b110010110100100111: begin rgb_reg = 3'b111; end
            18'b110010110100101010: begin rgb_reg = 3'b111; end
            18'b110010110100101011: begin rgb_reg = 3'b111; end
            18'b110010110100110010: begin rgb_reg = 3'b111; end
            18'b110010110100110011: begin rgb_reg = 3'b111; end
            18'b110010110100111000: begin rgb_reg = 3'b111; end
            18'b110010110100111001: begin rgb_reg = 3'b111; end
            18'b110010110100111010: begin rgb_reg = 3'b111; end
            18'b110010110100111011: begin rgb_reg = 3'b111; end
            18'b110010110100111100: begin rgb_reg = 3'b111; end
            18'b110010110100111101: begin rgb_reg = 3'b111; end
            18'b110010110100111110: begin rgb_reg = 3'b111; end
            18'b110010110100111111: begin rgb_reg = 3'b111; end
            18'b110010110101000010: begin rgb_reg = 3'b111; end
            18'b110010110101000011: begin rgb_reg = 3'b111; end
            18'b110010110101001010: begin rgb_reg = 3'b111; end
            18'b110010110101001011: begin rgb_reg = 3'b111; end
            18'b110010110101001110: begin rgb_reg = 3'b111; end
            18'b110010110101001111: begin rgb_reg = 3'b111; end
            18'b110010110101010010: begin rgb_reg = 3'b111; end
            18'b110010110101010011: begin rgb_reg = 3'b111; end
            18'b110010110101011110: begin rgb_reg = 3'b111; end
            18'b110010110101011111: begin rgb_reg = 3'b111; end
            18'b110010110101100110: begin rgb_reg = 3'b111; end
            18'b110010110101100111: begin rgb_reg = 3'b111; end
            18'b110010111010011000: begin rgb_reg = 3'b111; end
            18'b110010111010011001: begin rgb_reg = 3'b111; end
            18'b110010111010100000: begin rgb_reg = 3'b111; end
            18'b110010111010100001: begin rgb_reg = 3'b111; end
            18'b110010111010100110: begin rgb_reg = 3'b111; end
            18'b110010111010100111: begin rgb_reg = 3'b111; end
            18'b110010111010101000: begin rgb_reg = 3'b111; end
            18'b110010111010101001: begin rgb_reg = 3'b111; end
            18'b110010111010101010: begin rgb_reg = 3'b111; end
            18'b110010111010101011: begin rgb_reg = 3'b111; end
            18'b110010111010101100: begin rgb_reg = 3'b111; end
            18'b110010111010101101: begin rgb_reg = 3'b111; end
            18'b110010111010110000: begin rgb_reg = 3'b111; end
            18'b110010111010110001: begin rgb_reg = 3'b111; end
            18'b110010111010111100: begin rgb_reg = 3'b111; end
            18'b110010111010111101: begin rgb_reg = 3'b111; end
            18'b110010111011000000: begin rgb_reg = 3'b111; end
            18'b110010111011000001: begin rgb_reg = 3'b111; end
            18'b110010111011001000: begin rgb_reg = 3'b111; end
            18'b110010111011001001: begin rgb_reg = 3'b111; end
            18'b110010111011011100: begin rgb_reg = 3'b111; end
            18'b110010111011011101: begin rgb_reg = 3'b111; end
            18'b110010111011100100: begin rgb_reg = 3'b111; end
            18'b110010111011100101: begin rgb_reg = 3'b111; end
            18'b110010111011110010: begin rgb_reg = 3'b111; end
            18'b110010111011110011: begin rgb_reg = 3'b111; end
            18'b110010111011110100: begin rgb_reg = 3'b111; end
            18'b110010111011110101: begin rgb_reg = 3'b111; end
            18'b110010111011110110: begin rgb_reg = 3'b111; end
            18'b110010111011110111: begin rgb_reg = 3'b111; end
            18'b110010111011111000: begin rgb_reg = 3'b111; end
            18'b110010111011111001: begin rgb_reg = 3'b111; end
            18'b110010111011111100: begin rgb_reg = 3'b111; end
            18'b110010111011111101: begin rgb_reg = 3'b111; end
            18'b110010111011111110: begin rgb_reg = 3'b111; end
            18'b110010111011111111: begin rgb_reg = 3'b111; end
            18'b110010111100001000: begin rgb_reg = 3'b111; end
            18'b110010111100001001: begin rgb_reg = 3'b111; end
            18'b110010111100001010: begin rgb_reg = 3'b111; end
            18'b110010111100001011: begin rgb_reg = 3'b111; end
            18'b110010111100001100: begin rgb_reg = 3'b111; end
            18'b110010111100001101: begin rgb_reg = 3'b111; end
            18'b110010111100001110: begin rgb_reg = 3'b111; end
            18'b110010111100001111: begin rgb_reg = 3'b111; end
            18'b110010111100010010: begin rgb_reg = 3'b111; end
            18'b110010111100010011: begin rgb_reg = 3'b111; end
            18'b110010111100011110: begin rgb_reg = 3'b111; end
            18'b110010111100011111: begin rgb_reg = 3'b111; end
            18'b110010111100100110: begin rgb_reg = 3'b111; end
            18'b110010111100100111: begin rgb_reg = 3'b111; end
            18'b110010111100101010: begin rgb_reg = 3'b111; end
            18'b110010111100101011: begin rgb_reg = 3'b111; end
            18'b110010111100110010: begin rgb_reg = 3'b111; end
            18'b110010111100110011: begin rgb_reg = 3'b111; end
            18'b110010111100111000: begin rgb_reg = 3'b111; end
            18'b110010111100111001: begin rgb_reg = 3'b111; end
            18'b110010111100111010: begin rgb_reg = 3'b111; end
            18'b110010111100111011: begin rgb_reg = 3'b111; end
            18'b110010111100111100: begin rgb_reg = 3'b111; end
            18'b110010111100111101: begin rgb_reg = 3'b111; end
            18'b110010111100111110: begin rgb_reg = 3'b111; end
            18'b110010111100111111: begin rgb_reg = 3'b111; end
            18'b110010111101000010: begin rgb_reg = 3'b111; end
            18'b110010111101000011: begin rgb_reg = 3'b111; end
            18'b110010111101001010: begin rgb_reg = 3'b111; end
            18'b110010111101001011: begin rgb_reg = 3'b111; end
            18'b110010111101001110: begin rgb_reg = 3'b111; end
            18'b110010111101001111: begin rgb_reg = 3'b111; end
            18'b110010111101010010: begin rgb_reg = 3'b111; end
            18'b110010111101010011: begin rgb_reg = 3'b111; end
            18'b110010111101011110: begin rgb_reg = 3'b111; end
            18'b110010111101011111: begin rgb_reg = 3'b111; end
            18'b110010111101100110: begin rgb_reg = 3'b111; end
            18'b110010111101100111: begin rgb_reg = 3'b111; end
            18'b110011000010011000: begin rgb_reg = 3'b111; end
            18'b110011000010011001: begin rgb_reg = 3'b111; end
            18'b110011000010100000: begin rgb_reg = 3'b111; end
            18'b110011000010100001: begin rgb_reg = 3'b111; end
            18'b110011000010100100: begin rgb_reg = 3'b111; end
            18'b110011000010100101: begin rgb_reg = 3'b111; end
            18'b110011000010101100: begin rgb_reg = 3'b111; end
            18'b110011000010101101: begin rgb_reg = 3'b111; end
            18'b110011000010110000: begin rgb_reg = 3'b111; end
            18'b110011000010110001: begin rgb_reg = 3'b111; end
            18'b110011000010111100: begin rgb_reg = 3'b111; end
            18'b110011000010111101: begin rgb_reg = 3'b111; end
            18'b110011000011000000: begin rgb_reg = 3'b111; end
            18'b110011000011000001: begin rgb_reg = 3'b111; end
            18'b110011000011001000: begin rgb_reg = 3'b111; end
            18'b110011000011001001: begin rgb_reg = 3'b111; end
            18'b110011000011011100: begin rgb_reg = 3'b111; end
            18'b110011000011011101: begin rgb_reg = 3'b111; end
            18'b110011000011100100: begin rgb_reg = 3'b111; end
            18'b110011000011100101: begin rgb_reg = 3'b111; end
            18'b110011000011110000: begin rgb_reg = 3'b111; end
            18'b110011000011110001: begin rgb_reg = 3'b111; end
            18'b110011000011111000: begin rgb_reg = 3'b111; end
            18'b110011000011111001: begin rgb_reg = 3'b111; end
            18'b110011000011111100: begin rgb_reg = 3'b111; end
            18'b110011000011111101: begin rgb_reg = 3'b111; end
            18'b110011000100000000: begin rgb_reg = 3'b111; end
            18'b110011000100000001: begin rgb_reg = 3'b111; end
            18'b110011000100000110: begin rgb_reg = 3'b111; end
            18'b110011000100000111: begin rgb_reg = 3'b111; end
            18'b110011000100001110: begin rgb_reg = 3'b111; end
            18'b110011000100001111: begin rgb_reg = 3'b111; end
            18'b110011000100010010: begin rgb_reg = 3'b111; end
            18'b110011000100010011: begin rgb_reg = 3'b111; end
            18'b110011000100011110: begin rgb_reg = 3'b111; end
            18'b110011000100011111: begin rgb_reg = 3'b111; end
            18'b110011000100100110: begin rgb_reg = 3'b111; end
            18'b110011000100100111: begin rgb_reg = 3'b111; end
            18'b110011000100101100: begin rgb_reg = 3'b111; end
            18'b110011000100101101: begin rgb_reg = 3'b111; end
            18'b110011000100110000: begin rgb_reg = 3'b111; end
            18'b110011000100110001: begin rgb_reg = 3'b111; end
            18'b110011000100110110: begin rgb_reg = 3'b111; end
            18'b110011000100110111: begin rgb_reg = 3'b111; end
            18'b110011000100111110: begin rgb_reg = 3'b111; end
            18'b110011000100111111: begin rgb_reg = 3'b111; end
            18'b110011000101000010: begin rgb_reg = 3'b111; end
            18'b110011000101000011: begin rgb_reg = 3'b111; end
            18'b110011000101001010: begin rgb_reg = 3'b111; end
            18'b110011000101001011: begin rgb_reg = 3'b111; end
            18'b110011000101001110: begin rgb_reg = 3'b111; end
            18'b110011000101001111: begin rgb_reg = 3'b111; end
            18'b110011000101010010: begin rgb_reg = 3'b111; end
            18'b110011000101010011: begin rgb_reg = 3'b111; end
            18'b110011000101011010: begin rgb_reg = 3'b111; end
            18'b110011000101011011: begin rgb_reg = 3'b111; end
            18'b110011000101011110: begin rgb_reg = 3'b111; end
            18'b110011000101011111: begin rgb_reg = 3'b111; end
            18'b110011000101100110: begin rgb_reg = 3'b111; end
            18'b110011000101100111: begin rgb_reg = 3'b111; end
            18'b110011001010011000: begin rgb_reg = 3'b111; end
            18'b110011001010011001: begin rgb_reg = 3'b111; end
            18'b110011001010100000: begin rgb_reg = 3'b111; end
            18'b110011001010100001: begin rgb_reg = 3'b111; end
            18'b110011001010100100: begin rgb_reg = 3'b111; end
            18'b110011001010100101: begin rgb_reg = 3'b111; end
            18'b110011001010101100: begin rgb_reg = 3'b111; end
            18'b110011001010101101: begin rgb_reg = 3'b111; end
            18'b110011001010110000: begin rgb_reg = 3'b111; end
            18'b110011001010110001: begin rgb_reg = 3'b111; end
            18'b110011001010111100: begin rgb_reg = 3'b111; end
            18'b110011001010111101: begin rgb_reg = 3'b111; end
            18'b110011001011000000: begin rgb_reg = 3'b111; end
            18'b110011001011000001: begin rgb_reg = 3'b111; end
            18'b110011001011001000: begin rgb_reg = 3'b111; end
            18'b110011001011001001: begin rgb_reg = 3'b111; end
            18'b110011001011011100: begin rgb_reg = 3'b111; end
            18'b110011001011011101: begin rgb_reg = 3'b111; end
            18'b110011001011100100: begin rgb_reg = 3'b111; end
            18'b110011001011100101: begin rgb_reg = 3'b111; end
            18'b110011001011110000: begin rgb_reg = 3'b111; end
            18'b110011001011110001: begin rgb_reg = 3'b111; end
            18'b110011001011111000: begin rgb_reg = 3'b111; end
            18'b110011001011111001: begin rgb_reg = 3'b111; end
            18'b110011001011111100: begin rgb_reg = 3'b111; end
            18'b110011001011111101: begin rgb_reg = 3'b111; end
            18'b110011001100000000: begin rgb_reg = 3'b111; end
            18'b110011001100000001: begin rgb_reg = 3'b111; end
            18'b110011001100000110: begin rgb_reg = 3'b111; end
            18'b110011001100000111: begin rgb_reg = 3'b111; end
            18'b110011001100001110: begin rgb_reg = 3'b111; end
            18'b110011001100001111: begin rgb_reg = 3'b111; end
            18'b110011001100010010: begin rgb_reg = 3'b111; end
            18'b110011001100010011: begin rgb_reg = 3'b111; end
            18'b110011001100011110: begin rgb_reg = 3'b111; end
            18'b110011001100011111: begin rgb_reg = 3'b111; end
            18'b110011001100100110: begin rgb_reg = 3'b111; end
            18'b110011001100100111: begin rgb_reg = 3'b111; end
            18'b110011001100101100: begin rgb_reg = 3'b111; end
            18'b110011001100101101: begin rgb_reg = 3'b111; end
            18'b110011001100110000: begin rgb_reg = 3'b111; end
            18'b110011001100110001: begin rgb_reg = 3'b111; end
            18'b110011001100110110: begin rgb_reg = 3'b111; end
            18'b110011001100110111: begin rgb_reg = 3'b111; end
            18'b110011001100111110: begin rgb_reg = 3'b111; end
            18'b110011001100111111: begin rgb_reg = 3'b111; end
            18'b110011001101000010: begin rgb_reg = 3'b111; end
            18'b110011001101000011: begin rgb_reg = 3'b111; end
            18'b110011001101001010: begin rgb_reg = 3'b111; end
            18'b110011001101001011: begin rgb_reg = 3'b111; end
            18'b110011001101001110: begin rgb_reg = 3'b111; end
            18'b110011001101001111: begin rgb_reg = 3'b111; end
            18'b110011001101010010: begin rgb_reg = 3'b111; end
            18'b110011001101010011: begin rgb_reg = 3'b111; end
            18'b110011001101011010: begin rgb_reg = 3'b111; end
            18'b110011001101011011: begin rgb_reg = 3'b111; end
            18'b110011001101011110: begin rgb_reg = 3'b111; end
            18'b110011001101011111: begin rgb_reg = 3'b111; end
            18'b110011001101100110: begin rgb_reg = 3'b111; end
            18'b110011001101100111: begin rgb_reg = 3'b111; end
            18'b110011010010011000: begin rgb_reg = 3'b111; end
            18'b110011010010011001: begin rgb_reg = 3'b111; end
            18'b110011010010100000: begin rgb_reg = 3'b111; end
            18'b110011010010100001: begin rgb_reg = 3'b111; end
            18'b110011010010100110: begin rgb_reg = 3'b111; end
            18'b110011010010100111: begin rgb_reg = 3'b111; end
            18'b110011010010101000: begin rgb_reg = 3'b111; end
            18'b110011010010101001: begin rgb_reg = 3'b111; end
            18'b110011010010101010: begin rgb_reg = 3'b111; end
            18'b110011010010101011: begin rgb_reg = 3'b111; end
            18'b110011010010101100: begin rgb_reg = 3'b111; end
            18'b110011010010101101: begin rgb_reg = 3'b111; end
            18'b110011010010110000: begin rgb_reg = 3'b111; end
            18'b110011010010110001: begin rgb_reg = 3'b111; end
            18'b110011010010111100: begin rgb_reg = 3'b111; end
            18'b110011010010111101: begin rgb_reg = 3'b111; end
            18'b110011010011000000: begin rgb_reg = 3'b111; end
            18'b110011010011000001: begin rgb_reg = 3'b111; end
            18'b110011010011001000: begin rgb_reg = 3'b111; end
            18'b110011010011001001: begin rgb_reg = 3'b111; end
            18'b110011010011011100: begin rgb_reg = 3'b111; end
            18'b110011010011011101: begin rgb_reg = 3'b111; end
            18'b110011010011100100: begin rgb_reg = 3'b111; end
            18'b110011010011100101: begin rgb_reg = 3'b111; end
            18'b110011010011110010: begin rgb_reg = 3'b111; end
            18'b110011010011110011: begin rgb_reg = 3'b111; end
            18'b110011010011110100: begin rgb_reg = 3'b111; end
            18'b110011010011110101: begin rgb_reg = 3'b111; end
            18'b110011010011110110: begin rgb_reg = 3'b111; end
            18'b110011010011110111: begin rgb_reg = 3'b111; end
            18'b110011010011111000: begin rgb_reg = 3'b111; end
            18'b110011010011111001: begin rgb_reg = 3'b111; end
            18'b110011010011111100: begin rgb_reg = 3'b111; end
            18'b110011010011111101: begin rgb_reg = 3'b111; end
            18'b110011010100000010: begin rgb_reg = 3'b111; end
            18'b110011010100000011: begin rgb_reg = 3'b111; end
            18'b110011010100001000: begin rgb_reg = 3'b111; end
            18'b110011010100001001: begin rgb_reg = 3'b111; end
            18'b110011010100001010: begin rgb_reg = 3'b111; end
            18'b110011010100001011: begin rgb_reg = 3'b111; end
            18'b110011010100001100: begin rgb_reg = 3'b111; end
            18'b110011010100001101: begin rgb_reg = 3'b111; end
            18'b110011010100001110: begin rgb_reg = 3'b111; end
            18'b110011010100001111: begin rgb_reg = 3'b111; end
            18'b110011010100010010: begin rgb_reg = 3'b111; end
            18'b110011010100010011: begin rgb_reg = 3'b111; end
            18'b110011010100011110: begin rgb_reg = 3'b111; end
            18'b110011010100011111: begin rgb_reg = 3'b111; end
            18'b110011010100100110: begin rgb_reg = 3'b111; end
            18'b110011010100100111: begin rgb_reg = 3'b111; end
            18'b110011010100101110: begin rgb_reg = 3'b111; end
            18'b110011010100101111: begin rgb_reg = 3'b111; end
            18'b110011010100111000: begin rgb_reg = 3'b111; end
            18'b110011010100111001: begin rgb_reg = 3'b111; end
            18'b110011010100111010: begin rgb_reg = 3'b111; end
            18'b110011010100111011: begin rgb_reg = 3'b111; end
            18'b110011010100111100: begin rgb_reg = 3'b111; end
            18'b110011010100111101: begin rgb_reg = 3'b111; end
            18'b110011010100111110: begin rgb_reg = 3'b111; end
            18'b110011010100111111: begin rgb_reg = 3'b111; end
            18'b110011010101000010: begin rgb_reg = 3'b111; end
            18'b110011010101000011: begin rgb_reg = 3'b111; end
            18'b110011010101001010: begin rgb_reg = 3'b111; end
            18'b110011010101001011: begin rgb_reg = 3'b111; end
            18'b110011010101001110: begin rgb_reg = 3'b111; end
            18'b110011010101001111: begin rgb_reg = 3'b111; end
            18'b110011010101010100: begin rgb_reg = 3'b111; end
            18'b110011010101010101: begin rgb_reg = 3'b111; end
            18'b110011010101010110: begin rgb_reg = 3'b111; end
            18'b110011010101010111: begin rgb_reg = 3'b111; end
            18'b110011010101011000: begin rgb_reg = 3'b111; end
            18'b110011010101011001: begin rgb_reg = 3'b111; end
            18'b110011010101011110: begin rgb_reg = 3'b111; end
            18'b110011010101011111: begin rgb_reg = 3'b111; end
            18'b110011010101100110: begin rgb_reg = 3'b111; end
            18'b110011010101100111: begin rgb_reg = 3'b111; end
            18'b110011011010011000: begin rgb_reg = 3'b111; end
            18'b110011011010011001: begin rgb_reg = 3'b111; end
            18'b110011011010100000: begin rgb_reg = 3'b111; end
            18'b110011011010100001: begin rgb_reg = 3'b111; end
            18'b110011011010100110: begin rgb_reg = 3'b111; end
            18'b110011011010100111: begin rgb_reg = 3'b111; end
            18'b110011011010101000: begin rgb_reg = 3'b111; end
            18'b110011011010101001: begin rgb_reg = 3'b111; end
            18'b110011011010101010: begin rgb_reg = 3'b111; end
            18'b110011011010101011: begin rgb_reg = 3'b111; end
            18'b110011011010101100: begin rgb_reg = 3'b111; end
            18'b110011011010101101: begin rgb_reg = 3'b111; end
            18'b110011011010110000: begin rgb_reg = 3'b111; end
            18'b110011011010110001: begin rgb_reg = 3'b111; end
            18'b110011011010111100: begin rgb_reg = 3'b111; end
            18'b110011011010111101: begin rgb_reg = 3'b111; end
            18'b110011011011000000: begin rgb_reg = 3'b111; end
            18'b110011011011000001: begin rgb_reg = 3'b111; end
            18'b110011011011001000: begin rgb_reg = 3'b111; end
            18'b110011011011001001: begin rgb_reg = 3'b111; end
            18'b110011011011011100: begin rgb_reg = 3'b111; end
            18'b110011011011011101: begin rgb_reg = 3'b111; end
            18'b110011011011100100: begin rgb_reg = 3'b111; end
            18'b110011011011100101: begin rgb_reg = 3'b111; end
            18'b110011011011110010: begin rgb_reg = 3'b111; end
            18'b110011011011110011: begin rgb_reg = 3'b111; end
            18'b110011011011110100: begin rgb_reg = 3'b111; end
            18'b110011011011110101: begin rgb_reg = 3'b111; end
            18'b110011011011110110: begin rgb_reg = 3'b111; end
            18'b110011011011110111: begin rgb_reg = 3'b111; end
            18'b110011011011111000: begin rgb_reg = 3'b111; end
            18'b110011011011111001: begin rgb_reg = 3'b111; end
            18'b110011011011111100: begin rgb_reg = 3'b111; end
            18'b110011011011111101: begin rgb_reg = 3'b111; end
            18'b110011011100000010: begin rgb_reg = 3'b111; end
            18'b110011011100000011: begin rgb_reg = 3'b111; end
            18'b110011011100001000: begin rgb_reg = 3'b111; end
            18'b110011011100001001: begin rgb_reg = 3'b111; end
            18'b110011011100001010: begin rgb_reg = 3'b111; end
            18'b110011011100001011: begin rgb_reg = 3'b111; end
            18'b110011011100001100: begin rgb_reg = 3'b111; end
            18'b110011011100001101: begin rgb_reg = 3'b111; end
            18'b110011011100001110: begin rgb_reg = 3'b111; end
            18'b110011011100001111: begin rgb_reg = 3'b111; end
            18'b110011011100010010: begin rgb_reg = 3'b111; end
            18'b110011011100010011: begin rgb_reg = 3'b111; end
            18'b110011011100011110: begin rgb_reg = 3'b111; end
            18'b110011011100011111: begin rgb_reg = 3'b111; end
            18'b110011011100100110: begin rgb_reg = 3'b111; end
            18'b110011011100100111: begin rgb_reg = 3'b111; end
            18'b110011011100101110: begin rgb_reg = 3'b111; end
            18'b110011011100101111: begin rgb_reg = 3'b111; end
            18'b110011011100111000: begin rgb_reg = 3'b111; end
            18'b110011011100111001: begin rgb_reg = 3'b111; end
            18'b110011011100111010: begin rgb_reg = 3'b111; end
            18'b110011011100111011: begin rgb_reg = 3'b111; end
            18'b110011011100111100: begin rgb_reg = 3'b111; end
            18'b110011011100111101: begin rgb_reg = 3'b111; end
            18'b110011011100111110: begin rgb_reg = 3'b111; end
            18'b110011011100111111: begin rgb_reg = 3'b111; end
            18'b110011011101000010: begin rgb_reg = 3'b111; end
            18'b110011011101000011: begin rgb_reg = 3'b111; end
            18'b110011011101001010: begin rgb_reg = 3'b111; end
            18'b110011011101001011: begin rgb_reg = 3'b111; end
            18'b110011011101001110: begin rgb_reg = 3'b111; end
            18'b110011011101001111: begin rgb_reg = 3'b111; end
            18'b110011011101010100: begin rgb_reg = 3'b111; end
            18'b110011011101010101: begin rgb_reg = 3'b111; end
            18'b110011011101010110: begin rgb_reg = 3'b111; end
            18'b110011011101010111: begin rgb_reg = 3'b111; end
            18'b110011011101011000: begin rgb_reg = 3'b111; end
            18'b110011011101011001: begin rgb_reg = 3'b111; end
            18'b110011011101011110: begin rgb_reg = 3'b111; end
            18'b110011011101011111: begin rgb_reg = 3'b111; end
            18'b110011011101100110: begin rgb_reg = 3'b111; end
            18'b110011011101100111: begin rgb_reg = 3'b111; end
            18'b110111100010010001: begin rgb_reg = 3'b101; end
            18'b110111100010010010: begin rgb_reg = 3'b101; end
            18'b110111100100001000: begin rgb_reg = 3'b101; end
            18'b110111100100001001: begin rgb_reg = 3'b101; end
            18'b110111101010010001: begin rgb_reg = 3'b101; end
            18'b110111101010010010: begin rgb_reg = 3'b101; end
            18'b110111101100001000: begin rgb_reg = 3'b101; end
            18'b110111101100001001: begin rgb_reg = 3'b101; end
            18'b110111110001101001: begin rgb_reg = 3'b101; end
            18'b110111110001101010: begin rgb_reg = 3'b101; end
            18'b110111110001110010: begin rgb_reg = 3'b101; end
            18'b110111110001110011: begin rgb_reg = 3'b101; end
            18'b110111110001110110: begin rgb_reg = 3'b101; end
            18'b110111110001110111: begin rgb_reg = 3'b101; end
            18'b110111110001111000: begin rgb_reg = 3'b101; end
            18'b110111110001111001: begin rgb_reg = 3'b101; end
            18'b110111110001111010: begin rgb_reg = 3'b101; end
            18'b110111110001111011: begin rgb_reg = 3'b101; end
            18'b110111110001111100: begin rgb_reg = 3'b101; end
            18'b110111110001111111: begin rgb_reg = 3'b101; end
            18'b110111110010000000: begin rgb_reg = 3'b101; end
            18'b110111110010000001: begin rgb_reg = 3'b101; end
            18'b110111110010000010: begin rgb_reg = 3'b101; end
            18'b110111110010000011: begin rgb_reg = 3'b101; end
            18'b110111110010000100: begin rgb_reg = 3'b101; end
            18'b110111110010000101: begin rgb_reg = 3'b101; end
            18'b110111110010000110: begin rgb_reg = 3'b101; end
            18'b110111110010000111: begin rgb_reg = 3'b101; end
            18'b110111110010001000: begin rgb_reg = 3'b101; end
            18'b110111110010001001: begin rgb_reg = 3'b101; end
            18'b110111110010010011: begin rgb_reg = 3'b101; end
            18'b110111110010010100: begin rgb_reg = 3'b101; end
            18'b110111110010011010: begin rgb_reg = 3'b101; end
            18'b110111110010011011: begin rgb_reg = 3'b101; end
            18'b110111110010011100: begin rgb_reg = 3'b101; end
            18'b110111110010011101: begin rgb_reg = 3'b101; end
            18'b110111110010011110: begin rgb_reg = 3'b101; end
            18'b110111110010011111: begin rgb_reg = 3'b101; end
            18'b110111110010100000: begin rgb_reg = 3'b101; end
            18'b110111110010100001: begin rgb_reg = 3'b101; end
            18'b110111110010100010: begin rgb_reg = 3'b101; end
            18'b110111110010100101: begin rgb_reg = 3'b101; end
            18'b110111110010100110: begin rgb_reg = 3'b101; end
            18'b110111110010100111: begin rgb_reg = 3'b101; end
            18'b110111110010101000: begin rgb_reg = 3'b101; end
            18'b110111110010101001: begin rgb_reg = 3'b101; end
            18'b110111110010101010: begin rgb_reg = 3'b101; end
            18'b110111110010101011: begin rgb_reg = 3'b101; end
            18'b110111110010101100: begin rgb_reg = 3'b101; end
            18'b110111110010101101: begin rgb_reg = 3'b101; end
            18'b110111110010110101: begin rgb_reg = 3'b101; end
            18'b110111110010110110: begin rgb_reg = 3'b101; end
            18'b110111110010110111: begin rgb_reg = 3'b101; end
            18'b110111110010111000: begin rgb_reg = 3'b101; end
            18'b110111110010111001: begin rgb_reg = 3'b101; end
            18'b110111110010111010: begin rgb_reg = 3'b101; end
            18'b110111110010111011: begin rgb_reg = 3'b101; end
            18'b110111110011000011: begin rgb_reg = 3'b101; end
            18'b110111110011000100: begin rgb_reg = 3'b101; end
            18'b110111110011000101: begin rgb_reg = 3'b101; end
            18'b110111110011000110: begin rgb_reg = 3'b101; end
            18'b110111110011000111: begin rgb_reg = 3'b101; end
            18'b110111110011001000: begin rgb_reg = 3'b101; end
            18'b110111110011001110: begin rgb_reg = 3'b101; end
            18'b110111110011001111: begin rgb_reg = 3'b101; end
            18'b110111110011010000: begin rgb_reg = 3'b101; end
            18'b110111110011010001: begin rgb_reg = 3'b101; end
            18'b110111110011010010: begin rgb_reg = 3'b101; end
            18'b110111110011010011: begin rgb_reg = 3'b101; end
            18'b110111110011010100: begin rgb_reg = 3'b101; end
            18'b110111110011010101: begin rgb_reg = 3'b101; end
            18'b110111110011010110: begin rgb_reg = 3'b101; end
            18'b110111110011010111: begin rgb_reg = 3'b101; end
            18'b110111110011011000: begin rgb_reg = 3'b101; end
            18'b110111110011100000: begin rgb_reg = 3'b101; end
            18'b110111110011100001: begin rgb_reg = 3'b101; end
            18'b110111110011100010: begin rgb_reg = 3'b101; end
            18'b110111110011100011: begin rgb_reg = 3'b101; end
            18'b110111110011100100: begin rgb_reg = 3'b101; end
            18'b110111110011100101: begin rgb_reg = 3'b101; end
            18'b110111110011100110: begin rgb_reg = 3'b101; end
            18'b110111110011100111: begin rgb_reg = 3'b101; end
            18'b110111110011101000: begin rgb_reg = 3'b101; end
            18'b110111110011110000: begin rgb_reg = 3'b101; end
            18'b110111110011110001: begin rgb_reg = 3'b101; end
            18'b110111110011110010: begin rgb_reg = 3'b101; end
            18'b110111110011110011: begin rgb_reg = 3'b101; end
            18'b110111110011110100: begin rgb_reg = 3'b101; end
            18'b110111110011110101: begin rgb_reg = 3'b101; end
            18'b110111110011111011: begin rgb_reg = 3'b101; end
            18'b110111110011111100: begin rgb_reg = 3'b101; end
            18'b110111110011111101: begin rgb_reg = 3'b101; end
            18'b110111110011111110: begin rgb_reg = 3'b101; end
            18'b110111110011111111: begin rgb_reg = 3'b101; end
            18'b110111110100000000: begin rgb_reg = 3'b101; end
            18'b110111110100000001: begin rgb_reg = 3'b101; end
            18'b110111110100000010: begin rgb_reg = 3'b101; end
            18'b110111110100000011: begin rgb_reg = 3'b101; end
            18'b110111110100001011: begin rgb_reg = 3'b101; end
            18'b110111110100001100: begin rgb_reg = 3'b101; end
            18'b110111110100010100: begin rgb_reg = 3'b101; end
            18'b110111110100010101: begin rgb_reg = 3'b101; end
            18'b110111110100010110: begin rgb_reg = 3'b101; end
            18'b110111110100010111: begin rgb_reg = 3'b101; end
            18'b110111110100011000: begin rgb_reg = 3'b101; end
            18'b110111110100011001: begin rgb_reg = 3'b101; end
            18'b110111110100011010: begin rgb_reg = 3'b101; end
            18'b110111110100011011: begin rgb_reg = 3'b101; end
            18'b110111110100011100: begin rgb_reg = 3'b101; end
            18'b110111110100011101: begin rgb_reg = 3'b101; end
            18'b110111110100011110: begin rgb_reg = 3'b101; end
            18'b110111110100100011: begin rgb_reg = 3'b101; end
            18'b110111110100100100: begin rgb_reg = 3'b101; end
            18'b110111110100100101: begin rgb_reg = 3'b101; end
            18'b110111110100100110: begin rgb_reg = 3'b101; end
            18'b110111110100100111: begin rgb_reg = 3'b101; end
            18'b110111110100101000: begin rgb_reg = 3'b101; end
            18'b110111110100101001: begin rgb_reg = 3'b101; end
            18'b110111110100110101: begin rgb_reg = 3'b101; end
            18'b110111110100110110: begin rgb_reg = 3'b101; end
            18'b110111110100110111: begin rgb_reg = 3'b101; end
            18'b110111110100111000: begin rgb_reg = 3'b101; end
            18'b110111110100111001: begin rgb_reg = 3'b101; end
            18'b110111110100111010: begin rgb_reg = 3'b101; end
            18'b110111110100111011: begin rgb_reg = 3'b101; end
            18'b110111110101000011: begin rgb_reg = 3'b101; end
            18'b110111110101000100: begin rgb_reg = 3'b101; end
            18'b110111110101000101: begin rgb_reg = 3'b101; end
            18'b110111110101000110: begin rgb_reg = 3'b101; end
            18'b110111110101000111: begin rgb_reg = 3'b101; end
            18'b110111110101001000: begin rgb_reg = 3'b101; end
            18'b110111110101001110: begin rgb_reg = 3'b101; end
            18'b110111110101001111: begin rgb_reg = 3'b101; end
            18'b110111110101010111: begin rgb_reg = 3'b101; end
            18'b110111110101011000: begin rgb_reg = 3'b101; end
            18'b110111110101011100: begin rgb_reg = 3'b101; end
            18'b110111110101011101: begin rgb_reg = 3'b101; end
            18'b110111110101011110: begin rgb_reg = 3'b101; end
            18'b110111110101011111: begin rgb_reg = 3'b101; end
            18'b110111110101100000: begin rgb_reg = 3'b101; end
            18'b110111110101100001: begin rgb_reg = 3'b101; end
            18'b110111110101100010: begin rgb_reg = 3'b101; end
            18'b110111110101100011: begin rgb_reg = 3'b101; end
            18'b110111110101100100: begin rgb_reg = 3'b101; end
            18'b110111110101100101: begin rgb_reg = 3'b101; end
            18'b110111110101100110: begin rgb_reg = 3'b101; end
            18'b110111110101101001: begin rgb_reg = 3'b101; end
            18'b110111110101101010: begin rgb_reg = 3'b101; end
            18'b110111110101101011: begin rgb_reg = 3'b101; end
            18'b110111110101101100: begin rgb_reg = 3'b101; end
            18'b110111110101101101: begin rgb_reg = 3'b101; end
            18'b110111110101101110: begin rgb_reg = 3'b101; end
            18'b110111110101101111: begin rgb_reg = 3'b101; end
            18'b110111110101110010: begin rgb_reg = 3'b101; end
            18'b110111110101110011: begin rgb_reg = 3'b101; end
            18'b110111110101111011: begin rgb_reg = 3'b101; end
            18'b110111110101111100: begin rgb_reg = 3'b101; end
            18'b110111110110000000: begin rgb_reg = 3'b101; end
            18'b110111110110000001: begin rgb_reg = 3'b101; end
            18'b110111110110001001: begin rgb_reg = 3'b101; end
            18'b110111110110001010: begin rgb_reg = 3'b101; end
            18'b110111110110001101: begin rgb_reg = 3'b101; end
            18'b110111110110001110: begin rgb_reg = 3'b101; end
            18'b110111110110001111: begin rgb_reg = 3'b101; end
            18'b110111110110010000: begin rgb_reg = 3'b101; end
            18'b110111110110010001: begin rgb_reg = 3'b101; end
            18'b110111110110010010: begin rgb_reg = 3'b101; end
            18'b110111110110010011: begin rgb_reg = 3'b101; end
            18'b110111110110010100: begin rgb_reg = 3'b101; end
            18'b110111110110010101: begin rgb_reg = 3'b101; end
            18'b110111110110010110: begin rgb_reg = 3'b101; end
            18'b110111110110010111: begin rgb_reg = 3'b101; end
            18'b110111111001101001: begin rgb_reg = 3'b101; end
            18'b110111111001101010: begin rgb_reg = 3'b101; end
            18'b110111111001110010: begin rgb_reg = 3'b101; end
            18'b110111111001110011: begin rgb_reg = 3'b101; end
            18'b110111111001110110: begin rgb_reg = 3'b101; end
            18'b110111111001110111: begin rgb_reg = 3'b101; end
            18'b110111111001111000: begin rgb_reg = 3'b101; end
            18'b110111111001111001: begin rgb_reg = 3'b101; end
            18'b110111111001111010: begin rgb_reg = 3'b101; end
            18'b110111111001111011: begin rgb_reg = 3'b101; end
            18'b110111111001111100: begin rgb_reg = 3'b101; end
            18'b110111111001111111: begin rgb_reg = 3'b101; end
            18'b110111111010000000: begin rgb_reg = 3'b101; end
            18'b110111111010000001: begin rgb_reg = 3'b101; end
            18'b110111111010000010: begin rgb_reg = 3'b101; end
            18'b110111111010000011: begin rgb_reg = 3'b101; end
            18'b110111111010000100: begin rgb_reg = 3'b101; end
            18'b110111111010000101: begin rgb_reg = 3'b101; end
            18'b110111111010000110: begin rgb_reg = 3'b101; end
            18'b110111111010000111: begin rgb_reg = 3'b101; end
            18'b110111111010001000: begin rgb_reg = 3'b101; end
            18'b110111111010001001: begin rgb_reg = 3'b101; end
            18'b110111111010010011: begin rgb_reg = 3'b101; end
            18'b110111111010010100: begin rgb_reg = 3'b101; end
            18'b110111111010011010: begin rgb_reg = 3'b101; end
            18'b110111111010011011: begin rgb_reg = 3'b101; end
            18'b110111111010011100: begin rgb_reg = 3'b101; end
            18'b110111111010011101: begin rgb_reg = 3'b101; end
            18'b110111111010011110: begin rgb_reg = 3'b101; end
            18'b110111111010011111: begin rgb_reg = 3'b101; end
            18'b110111111010100000: begin rgb_reg = 3'b101; end
            18'b110111111010100001: begin rgb_reg = 3'b101; end
            18'b110111111010100010: begin rgb_reg = 3'b101; end
            18'b110111111010100101: begin rgb_reg = 3'b101; end
            18'b110111111010100110: begin rgb_reg = 3'b101; end
            18'b110111111010100111: begin rgb_reg = 3'b101; end
            18'b110111111010101000: begin rgb_reg = 3'b101; end
            18'b110111111010101001: begin rgb_reg = 3'b101; end
            18'b110111111010101010: begin rgb_reg = 3'b101; end
            18'b110111111010101011: begin rgb_reg = 3'b101; end
            18'b110111111010101100: begin rgb_reg = 3'b101; end
            18'b110111111010101101: begin rgb_reg = 3'b101; end
            18'b110111111010110101: begin rgb_reg = 3'b101; end
            18'b110111111010110110: begin rgb_reg = 3'b101; end
            18'b110111111010110111: begin rgb_reg = 3'b101; end
            18'b110111111010111000: begin rgb_reg = 3'b101; end
            18'b110111111010111001: begin rgb_reg = 3'b101; end
            18'b110111111010111010: begin rgb_reg = 3'b101; end
            18'b110111111010111011: begin rgb_reg = 3'b101; end
            18'b110111111011000011: begin rgb_reg = 3'b101; end
            18'b110111111011000100: begin rgb_reg = 3'b101; end
            18'b110111111011000101: begin rgb_reg = 3'b101; end
            18'b110111111011000110: begin rgb_reg = 3'b101; end
            18'b110111111011000111: begin rgb_reg = 3'b101; end
            18'b110111111011001000: begin rgb_reg = 3'b101; end
            18'b110111111011001110: begin rgb_reg = 3'b101; end
            18'b110111111011001111: begin rgb_reg = 3'b101; end
            18'b110111111011010000: begin rgb_reg = 3'b101; end
            18'b110111111011010001: begin rgb_reg = 3'b101; end
            18'b110111111011010010: begin rgb_reg = 3'b101; end
            18'b110111111011010011: begin rgb_reg = 3'b101; end
            18'b110111111011010100: begin rgb_reg = 3'b101; end
            18'b110111111011010101: begin rgb_reg = 3'b101; end
            18'b110111111011010110: begin rgb_reg = 3'b101; end
            18'b110111111011010111: begin rgb_reg = 3'b101; end
            18'b110111111011011000: begin rgb_reg = 3'b101; end
            18'b110111111011100000: begin rgb_reg = 3'b101; end
            18'b110111111011100001: begin rgb_reg = 3'b101; end
            18'b110111111011100010: begin rgb_reg = 3'b101; end
            18'b110111111011100011: begin rgb_reg = 3'b101; end
            18'b110111111011100100: begin rgb_reg = 3'b101; end
            18'b110111111011100101: begin rgb_reg = 3'b101; end
            18'b110111111011100110: begin rgb_reg = 3'b101; end
            18'b110111111011100111: begin rgb_reg = 3'b101; end
            18'b110111111011101000: begin rgb_reg = 3'b101; end
            18'b110111111011110000: begin rgb_reg = 3'b101; end
            18'b110111111011110001: begin rgb_reg = 3'b101; end
            18'b110111111011110010: begin rgb_reg = 3'b101; end
            18'b110111111011110011: begin rgb_reg = 3'b101; end
            18'b110111111011110100: begin rgb_reg = 3'b101; end
            18'b110111111011110101: begin rgb_reg = 3'b101; end
            18'b110111111011111011: begin rgb_reg = 3'b101; end
            18'b110111111011111100: begin rgb_reg = 3'b101; end
            18'b110111111011111101: begin rgb_reg = 3'b101; end
            18'b110111111011111110: begin rgb_reg = 3'b101; end
            18'b110111111011111111: begin rgb_reg = 3'b101; end
            18'b110111111100000000: begin rgb_reg = 3'b101; end
            18'b110111111100000001: begin rgb_reg = 3'b101; end
            18'b110111111100000010: begin rgb_reg = 3'b101; end
            18'b110111111100000011: begin rgb_reg = 3'b101; end
            18'b110111111100001011: begin rgb_reg = 3'b101; end
            18'b110111111100001100: begin rgb_reg = 3'b101; end
            18'b110111111100010100: begin rgb_reg = 3'b101; end
            18'b110111111100010101: begin rgb_reg = 3'b101; end
            18'b110111111100010110: begin rgb_reg = 3'b101; end
            18'b110111111100010111: begin rgb_reg = 3'b101; end
            18'b110111111100011000: begin rgb_reg = 3'b101; end
            18'b110111111100011001: begin rgb_reg = 3'b101; end
            18'b110111111100011010: begin rgb_reg = 3'b101; end
            18'b110111111100011011: begin rgb_reg = 3'b101; end
            18'b110111111100011100: begin rgb_reg = 3'b101; end
            18'b110111111100011101: begin rgb_reg = 3'b101; end
            18'b110111111100011110: begin rgb_reg = 3'b101; end
            18'b110111111100100011: begin rgb_reg = 3'b101; end
            18'b110111111100100100: begin rgb_reg = 3'b101; end
            18'b110111111100100101: begin rgb_reg = 3'b101; end
            18'b110111111100100110: begin rgb_reg = 3'b101; end
            18'b110111111100100111: begin rgb_reg = 3'b101; end
            18'b110111111100101000: begin rgb_reg = 3'b101; end
            18'b110111111100101001: begin rgb_reg = 3'b101; end
            18'b110111111100110101: begin rgb_reg = 3'b101; end
            18'b110111111100110110: begin rgb_reg = 3'b101; end
            18'b110111111100110111: begin rgb_reg = 3'b101; end
            18'b110111111100111000: begin rgb_reg = 3'b101; end
            18'b110111111100111001: begin rgb_reg = 3'b101; end
            18'b110111111100111010: begin rgb_reg = 3'b101; end
            18'b110111111100111011: begin rgb_reg = 3'b101; end
            18'b110111111101000011: begin rgb_reg = 3'b101; end
            18'b110111111101000100: begin rgb_reg = 3'b101; end
            18'b110111111101000101: begin rgb_reg = 3'b101; end
            18'b110111111101000110: begin rgb_reg = 3'b101; end
            18'b110111111101000111: begin rgb_reg = 3'b101; end
            18'b110111111101001000: begin rgb_reg = 3'b101; end
            18'b110111111101001110: begin rgb_reg = 3'b101; end
            18'b110111111101001111: begin rgb_reg = 3'b101; end
            18'b110111111101010111: begin rgb_reg = 3'b101; end
            18'b110111111101011000: begin rgb_reg = 3'b101; end
            18'b110111111101011100: begin rgb_reg = 3'b101; end
            18'b110111111101011101: begin rgb_reg = 3'b101; end
            18'b110111111101011110: begin rgb_reg = 3'b101; end
            18'b110111111101011111: begin rgb_reg = 3'b101; end
            18'b110111111101100000: begin rgb_reg = 3'b101; end
            18'b110111111101100001: begin rgb_reg = 3'b101; end
            18'b110111111101100010: begin rgb_reg = 3'b101; end
            18'b110111111101100011: begin rgb_reg = 3'b101; end
            18'b110111111101100100: begin rgb_reg = 3'b101; end
            18'b110111111101100101: begin rgb_reg = 3'b101; end
            18'b110111111101100110: begin rgb_reg = 3'b101; end
            18'b110111111101101001: begin rgb_reg = 3'b101; end
            18'b110111111101101010: begin rgb_reg = 3'b101; end
            18'b110111111101101011: begin rgb_reg = 3'b101; end
            18'b110111111101101100: begin rgb_reg = 3'b101; end
            18'b110111111101101101: begin rgb_reg = 3'b101; end
            18'b110111111101101110: begin rgb_reg = 3'b101; end
            18'b110111111101101111: begin rgb_reg = 3'b101; end
            18'b110111111101110010: begin rgb_reg = 3'b101; end
            18'b110111111101110011: begin rgb_reg = 3'b101; end
            18'b110111111101111011: begin rgb_reg = 3'b101; end
            18'b110111111101111100: begin rgb_reg = 3'b101; end
            18'b110111111110000000: begin rgb_reg = 3'b101; end
            18'b110111111110000001: begin rgb_reg = 3'b101; end
            18'b110111111110001001: begin rgb_reg = 3'b101; end
            18'b110111111110001010: begin rgb_reg = 3'b101; end
            18'b110111111110001101: begin rgb_reg = 3'b101; end
            18'b110111111110001110: begin rgb_reg = 3'b101; end
            18'b110111111110001111: begin rgb_reg = 3'b101; end
            18'b110111111110010000: begin rgb_reg = 3'b101; end
            18'b110111111110010001: begin rgb_reg = 3'b101; end
            18'b110111111110010010: begin rgb_reg = 3'b101; end
            18'b110111111110010011: begin rgb_reg = 3'b101; end
            18'b110111111110010100: begin rgb_reg = 3'b101; end
            18'b110111111110010101: begin rgb_reg = 3'b101; end
            18'b110111111110010110: begin rgb_reg = 3'b101; end
            18'b110111111110010111: begin rgb_reg = 3'b101; end
            18'b111000000001101001: begin rgb_reg = 3'b101; end
            18'b111000000001101010: begin rgb_reg = 3'b101; end
            18'b111000000001110010: begin rgb_reg = 3'b101; end
            18'b111000000001110011: begin rgb_reg = 3'b101; end
            18'b111000000001111000: begin rgb_reg = 3'b101; end
            18'b111000000001111001: begin rgb_reg = 3'b101; end
            18'b111000000010000100: begin rgb_reg = 3'b101; end
            18'b111000000010000101: begin rgb_reg = 3'b101; end
            18'b111000000010011000: begin rgb_reg = 3'b101; end
            18'b111000000010011001: begin rgb_reg = 3'b101; end
            18'b111000000010100101: begin rgb_reg = 3'b101; end
            18'b111000000010100110: begin rgb_reg = 3'b101; end
            18'b111000000010101111: begin rgb_reg = 3'b101; end
            18'b111000000010110011: begin rgb_reg = 3'b101; end
            18'b111000000010110100: begin rgb_reg = 3'b101; end
            18'b111000000010111100: begin rgb_reg = 3'b101; end
            18'b111000000010111101: begin rgb_reg = 3'b101; end
            18'b111000000011000001: begin rgb_reg = 3'b101; end
            18'b111000000011001010: begin rgb_reg = 3'b101; end
            18'b111000000011001110: begin rgb_reg = 3'b101; end
            18'b111000000011001111: begin rgb_reg = 3'b101; end
            18'b111000000011100000: begin rgb_reg = 3'b101; end
            18'b111000000011100001: begin rgb_reg = 3'b101; end
            18'b111000000011101001: begin rgb_reg = 3'b101; end
            18'b111000000011101010: begin rgb_reg = 3'b101; end
            18'b111000000011101110: begin rgb_reg = 3'b101; end
            18'b111000000011110111: begin rgb_reg = 3'b101; end
            18'b111000000011111011: begin rgb_reg = 3'b101; end
            18'b111000000011111100: begin rgb_reg = 3'b101; end
            18'b111000000100000100: begin rgb_reg = 3'b101; end
            18'b111000000100000101: begin rgb_reg = 3'b101; end
            18'b111000000100011000: begin rgb_reg = 3'b101; end
            18'b111000000100011001: begin rgb_reg = 3'b101; end
            18'b111000000100100001: begin rgb_reg = 3'b101; end
            18'b111000000100100010: begin rgb_reg = 3'b101; end
            18'b111000000100101010: begin rgb_reg = 3'b101; end
            18'b111000000100101011: begin rgb_reg = 3'b101; end
            18'b111000000100110011: begin rgb_reg = 3'b101; end
            18'b111000000100110100: begin rgb_reg = 3'b101; end
            18'b111000000100111100: begin rgb_reg = 3'b101; end
            18'b111000000100111101: begin rgb_reg = 3'b101; end
            18'b111000000101000001: begin rgb_reg = 3'b101; end
            18'b111000000101001010: begin rgb_reg = 3'b101; end
            18'b111000000101001110: begin rgb_reg = 3'b101; end
            18'b111000000101001111: begin rgb_reg = 3'b101; end
            18'b111000000101010000: begin rgb_reg = 3'b101; end
            18'b111000000101010001: begin rgb_reg = 3'b101; end
            18'b111000000101010111: begin rgb_reg = 3'b101; end
            18'b111000000101011000: begin rgb_reg = 3'b101; end
            18'b111000000101100000: begin rgb_reg = 3'b101; end
            18'b111000000101100001: begin rgb_reg = 3'b101; end
            18'b111000000101101011: begin rgb_reg = 3'b101; end
            18'b111000000101101100: begin rgb_reg = 3'b101; end
            18'b111000000101110010: begin rgb_reg = 3'b101; end
            18'b111000000101110011: begin rgb_reg = 3'b101; end
            18'b111000000101110100: begin rgb_reg = 3'b101; end
            18'b111000000101110101: begin rgb_reg = 3'b101; end
            18'b111000000101111011: begin rgb_reg = 3'b101; end
            18'b111000000101111100: begin rgb_reg = 3'b101; end
            18'b111000000110000000: begin rgb_reg = 3'b101; end
            18'b111000000110000001: begin rgb_reg = 3'b101; end
            18'b111000000110001001: begin rgb_reg = 3'b101; end
            18'b111000000110001010: begin rgb_reg = 3'b101; end
            18'b111000000110001101: begin rgb_reg = 3'b101; end
            18'b111000000110001110: begin rgb_reg = 3'b101; end
            18'b111000001001101001: begin rgb_reg = 3'b101; end
            18'b111000001001101010: begin rgb_reg = 3'b101; end
            18'b111000001001110010: begin rgb_reg = 3'b101; end
            18'b111000001001110011: begin rgb_reg = 3'b101; end
            18'b111000001001111000: begin rgb_reg = 3'b101; end
            18'b111000001001111001: begin rgb_reg = 3'b101; end
            18'b111000001010000100: begin rgb_reg = 3'b101; end
            18'b111000001010000101: begin rgb_reg = 3'b101; end
            18'b111000001010011000: begin rgb_reg = 3'b101; end
            18'b111000001010011001: begin rgb_reg = 3'b101; end
            18'b111000001010100101: begin rgb_reg = 3'b101; end
            18'b111000001010100110: begin rgb_reg = 3'b101; end
            18'b111000001010101110: begin rgb_reg = 3'b101; end
            18'b111000001010101111: begin rgb_reg = 3'b101; end
            18'b111000001010110011: begin rgb_reg = 3'b101; end
            18'b111000001010110100: begin rgb_reg = 3'b101; end
            18'b111000001010111100: begin rgb_reg = 3'b101; end
            18'b111000001010111101: begin rgb_reg = 3'b101; end
            18'b111000001011000000: begin rgb_reg = 3'b101; end
            18'b111000001011000001: begin rgb_reg = 3'b101; end
            18'b111000001011001001: begin rgb_reg = 3'b101; end
            18'b111000001011001010: begin rgb_reg = 3'b101; end
            18'b111000001011001110: begin rgb_reg = 3'b101; end
            18'b111000001011001111: begin rgb_reg = 3'b101; end
            18'b111000001011100000: begin rgb_reg = 3'b101; end
            18'b111000001011100001: begin rgb_reg = 3'b101; end
            18'b111000001011101001: begin rgb_reg = 3'b101; end
            18'b111000001011101010: begin rgb_reg = 3'b101; end
            18'b111000001011101101: begin rgb_reg = 3'b101; end
            18'b111000001011101110: begin rgb_reg = 3'b101; end
            18'b111000001011110110: begin rgb_reg = 3'b101; end
            18'b111000001011110111: begin rgb_reg = 3'b101; end
            18'b111000001011111011: begin rgb_reg = 3'b101; end
            18'b111000001011111100: begin rgb_reg = 3'b101; end
            18'b111000001100000100: begin rgb_reg = 3'b101; end
            18'b111000001100000101: begin rgb_reg = 3'b101; end
            18'b111000001100011000: begin rgb_reg = 3'b101; end
            18'b111000001100011001: begin rgb_reg = 3'b101; end
            18'b111000001100100001: begin rgb_reg = 3'b101; end
            18'b111000001100100010: begin rgb_reg = 3'b101; end
            18'b111000001100101010: begin rgb_reg = 3'b101; end
            18'b111000001100101011: begin rgb_reg = 3'b101; end
            18'b111000001100110011: begin rgb_reg = 3'b101; end
            18'b111000001100110100: begin rgb_reg = 3'b101; end
            18'b111000001100111100: begin rgb_reg = 3'b101; end
            18'b111000001100111101: begin rgb_reg = 3'b101; end
            18'b111000001101000001: begin rgb_reg = 3'b101; end
            18'b111000001101000010: begin rgb_reg = 3'b101; end
            18'b111000001101001010: begin rgb_reg = 3'b101; end
            18'b111000001101001011: begin rgb_reg = 3'b101; end
            18'b111000001101001110: begin rgb_reg = 3'b101; end
            18'b111000001101001111: begin rgb_reg = 3'b101; end
            18'b111000001101010000: begin rgb_reg = 3'b101; end
            18'b111000001101010001: begin rgb_reg = 3'b101; end
            18'b111000001101010111: begin rgb_reg = 3'b101; end
            18'b111000001101011000: begin rgb_reg = 3'b101; end
            18'b111000001101100000: begin rgb_reg = 3'b101; end
            18'b111000001101100001: begin rgb_reg = 3'b101; end
            18'b111000001101101011: begin rgb_reg = 3'b101; end
            18'b111000001101101100: begin rgb_reg = 3'b101; end
            18'b111000001101110010: begin rgb_reg = 3'b101; end
            18'b111000001101110011: begin rgb_reg = 3'b101; end
            18'b111000001101110100: begin rgb_reg = 3'b101; end
            18'b111000001101110101: begin rgb_reg = 3'b101; end
            18'b111000001101111011: begin rgb_reg = 3'b101; end
            18'b111000001101111100: begin rgb_reg = 3'b101; end
            18'b111000001110000000: begin rgb_reg = 3'b101; end
            18'b111000001110000001: begin rgb_reg = 3'b101; end
            18'b111000001110001001: begin rgb_reg = 3'b101; end
            18'b111000001110001010: begin rgb_reg = 3'b101; end
            18'b111000001110001101: begin rgb_reg = 3'b101; end
            18'b111000001110001110: begin rgb_reg = 3'b101; end
            18'b111000010001101001: begin rgb_reg = 3'b101; end
            18'b111000010001101010: begin rgb_reg = 3'b101; end
            18'b111000010001110001: begin rgb_reg = 3'b101; end
            18'b111000010001110010: begin rgb_reg = 3'b101; end
            18'b111000010001110011: begin rgb_reg = 3'b101; end
            18'b111000010001111000: begin rgb_reg = 3'b101; end
            18'b111000010001111001: begin rgb_reg = 3'b101; end
            18'b111000010010000100: begin rgb_reg = 3'b101; end
            18'b111000010010000101: begin rgb_reg = 3'b101; end
            18'b111000010010100101: begin rgb_reg = 3'b101; end
            18'b111000010010100110: begin rgb_reg = 3'b101; end
            18'b111000010010100111: begin rgb_reg = 3'b101; end
            18'b111000010010110011: begin rgb_reg = 3'b101; end
            18'b111000010010110100: begin rgb_reg = 3'b101; end
            18'b111000010010111100: begin rgb_reg = 3'b101; end
            18'b111000010010111101: begin rgb_reg = 3'b101; end
            18'b111000010011000000: begin rgb_reg = 3'b101; end
            18'b111000010011000001: begin rgb_reg = 3'b101; end
            18'b111000010011001110: begin rgb_reg = 3'b101; end
            18'b111000010011001111: begin rgb_reg = 3'b101; end
            18'b111000010011100000: begin rgb_reg = 3'b101; end
            18'b111000010011100001: begin rgb_reg = 3'b101; end
            18'b111000010011101101: begin rgb_reg = 3'b101; end
            18'b111000010011101110: begin rgb_reg = 3'b101; end
            18'b111000010011101111: begin rgb_reg = 3'b101; end
            18'b111000010011110110: begin rgb_reg = 3'b101; end
            18'b111000010011110111: begin rgb_reg = 3'b101; end
            18'b111000010011111011: begin rgb_reg = 3'b101; end
            18'b111000010011111100: begin rgb_reg = 3'b101; end
            18'b111000010100011000: begin rgb_reg = 3'b101; end
            18'b111000010100011001: begin rgb_reg = 3'b101; end
            18'b111000010100100001: begin rgb_reg = 3'b101; end
            18'b111000010100100010: begin rgb_reg = 3'b101; end
            18'b111000010100101010: begin rgb_reg = 3'b101; end
            18'b111000010100101011: begin rgb_reg = 3'b101; end
            18'b111000010100110011: begin rgb_reg = 3'b101; end
            18'b111000010100110100: begin rgb_reg = 3'b101; end
            18'b111000010101000001: begin rgb_reg = 3'b101; end
            18'b111000010101000010: begin rgb_reg = 3'b101; end
            18'b111000010101001010: begin rgb_reg = 3'b101; end
            18'b111000010101001011: begin rgb_reg = 3'b101; end
            18'b111000010101001110: begin rgb_reg = 3'b101; end
            18'b111000010101001111: begin rgb_reg = 3'b101; end
            18'b111000010101010111: begin rgb_reg = 3'b101; end
            18'b111000010101011000: begin rgb_reg = 3'b101; end
            18'b111000010101100000: begin rgb_reg = 3'b101; end
            18'b111000010101100001: begin rgb_reg = 3'b101; end
            18'b111000010101101011: begin rgb_reg = 3'b101; end
            18'b111000010101101100: begin rgb_reg = 3'b101; end
            18'b111000010101110010: begin rgb_reg = 3'b101; end
            18'b111000010101110011: begin rgb_reg = 3'b101; end
            18'b111000010101111011: begin rgb_reg = 3'b101; end
            18'b111000010101111100: begin rgb_reg = 3'b101; end
            18'b111000010110000000: begin rgb_reg = 3'b101; end
            18'b111000010110000001: begin rgb_reg = 3'b101; end
            18'b111000010110001001: begin rgb_reg = 3'b101; end
            18'b111000010110001010: begin rgb_reg = 3'b101; end
            18'b111000010110001101: begin rgb_reg = 3'b101; end
            18'b111000010110001110: begin rgb_reg = 3'b101; end
            18'b111000011001101001: begin rgb_reg = 3'b101; end
            18'b111000011001101010: begin rgb_reg = 3'b101; end
            18'b111000011001101011: begin rgb_reg = 3'b101; end
            18'b111000011001101100: begin rgb_reg = 3'b101; end
            18'b111000011001101101: begin rgb_reg = 3'b101; end
            18'b111000011001101110: begin rgb_reg = 3'b101; end
            18'b111000011001101111: begin rgb_reg = 3'b101; end
            18'b111000011001110000: begin rgb_reg = 3'b101; end
            18'b111000011001110001: begin rgb_reg = 3'b101; end
            18'b111000011001110010: begin rgb_reg = 3'b101; end
            18'b111000011001110011: begin rgb_reg = 3'b101; end
            18'b111000011001111000: begin rgb_reg = 3'b101; end
            18'b111000011001111001: begin rgb_reg = 3'b101; end
            18'b111000011010000100: begin rgb_reg = 3'b101; end
            18'b111000011010000101: begin rgb_reg = 3'b101; end
            18'b111000011010011010: begin rgb_reg = 3'b101; end
            18'b111000011010011011: begin rgb_reg = 3'b101; end
            18'b111000011010011100: begin rgb_reg = 3'b101; end
            18'b111000011010011101: begin rgb_reg = 3'b101; end
            18'b111000011010011110: begin rgb_reg = 3'b101; end
            18'b111000011010011111: begin rgb_reg = 3'b101; end
            18'b111000011010100000: begin rgb_reg = 3'b101; end
            18'b111000011010100101: begin rgb_reg = 3'b101; end
            18'b111000011010100110: begin rgb_reg = 3'b101; end
            18'b111000011010100111: begin rgb_reg = 3'b101; end
            18'b111000011010101000: begin rgb_reg = 3'b101; end
            18'b111000011010101001: begin rgb_reg = 3'b101; end
            18'b111000011010101010: begin rgb_reg = 3'b101; end
            18'b111000011010101011: begin rgb_reg = 3'b101; end
            18'b111000011010101100: begin rgb_reg = 3'b101; end
            18'b111000011010101101: begin rgb_reg = 3'b101; end
            18'b111000011010110011: begin rgb_reg = 3'b101; end
            18'b111000011010110100: begin rgb_reg = 3'b101; end
            18'b111000011010110101: begin rgb_reg = 3'b101; end
            18'b111000011010110110: begin rgb_reg = 3'b101; end
            18'b111000011010110111: begin rgb_reg = 3'b101; end
            18'b111000011010111000: begin rgb_reg = 3'b101; end
            18'b111000011010111001: begin rgb_reg = 3'b101; end
            18'b111000011010111010: begin rgb_reg = 3'b101; end
            18'b111000011010111011: begin rgb_reg = 3'b101; end
            18'b111000011010111100: begin rgb_reg = 3'b101; end
            18'b111000011010111101: begin rgb_reg = 3'b101; end
            18'b111000011011000000: begin rgb_reg = 3'b101; end
            18'b111000011011000001: begin rgb_reg = 3'b101; end
            18'b111000011011001110: begin rgb_reg = 3'b101; end
            18'b111000011011001111: begin rgb_reg = 3'b101; end
            18'b111000011011010000: begin rgb_reg = 3'b101; end
            18'b111000011011010001: begin rgb_reg = 3'b101; end
            18'b111000011011010010: begin rgb_reg = 3'b101; end
            18'b111000011011010011: begin rgb_reg = 3'b101; end
            18'b111000011011100000: begin rgb_reg = 3'b101; end
            18'b111000011011100001: begin rgb_reg = 3'b101; end
            18'b111000011011100010: begin rgb_reg = 3'b101; end
            18'b111000011011100011: begin rgb_reg = 3'b101; end
            18'b111000011011100100: begin rgb_reg = 3'b101; end
            18'b111000011011100101: begin rgb_reg = 3'b101; end
            18'b111000011011100110: begin rgb_reg = 3'b101; end
            18'b111000011011100111: begin rgb_reg = 3'b101; end
            18'b111000011011101000: begin rgb_reg = 3'b101; end
            18'b111000011011101101: begin rgb_reg = 3'b101; end
            18'b111000011011101110: begin rgb_reg = 3'b101; end
            18'b111000011011101111: begin rgb_reg = 3'b101; end
            18'b111000011011110000: begin rgb_reg = 3'b101; end
            18'b111000011011110001: begin rgb_reg = 3'b101; end
            18'b111000011011110010: begin rgb_reg = 3'b101; end
            18'b111000011011110011: begin rgb_reg = 3'b101; end
            18'b111000011011110100: begin rgb_reg = 3'b101; end
            18'b111000011011110101: begin rgb_reg = 3'b101; end
            18'b111000011011110110: begin rgb_reg = 3'b101; end
            18'b111000011011110111: begin rgb_reg = 3'b101; end
            18'b111000011011111011: begin rgb_reg = 3'b101; end
            18'b111000011011111100: begin rgb_reg = 3'b101; end
            18'b111000011011111101: begin rgb_reg = 3'b101; end
            18'b111000011011111110: begin rgb_reg = 3'b101; end
            18'b111000011011111111: begin rgb_reg = 3'b101; end
            18'b111000011100000000: begin rgb_reg = 3'b101; end
            18'b111000011100000001: begin rgb_reg = 3'b101; end
            18'b111000011100000010: begin rgb_reg = 3'b101; end
            18'b111000011100000011: begin rgb_reg = 3'b101; end
            18'b111000011100011000: begin rgb_reg = 3'b101; end
            18'b111000011100011001: begin rgb_reg = 3'b101; end
            18'b111000011100100001: begin rgb_reg = 3'b101; end
            18'b111000011100100010: begin rgb_reg = 3'b101; end
            18'b111000011100101010: begin rgb_reg = 3'b101; end
            18'b111000011100101011: begin rgb_reg = 3'b101; end
            18'b111000011100110011: begin rgb_reg = 3'b101; end
            18'b111000011100110100: begin rgb_reg = 3'b101; end
            18'b111000011101000001: begin rgb_reg = 3'b101; end
            18'b111000011101000010: begin rgb_reg = 3'b101; end
            18'b111000011101001010: begin rgb_reg = 3'b101; end
            18'b111000011101001011: begin rgb_reg = 3'b101; end
            18'b111000011101001110: begin rgb_reg = 3'b101; end
            18'b111000011101001111: begin rgb_reg = 3'b101; end
            18'b111000011101010011: begin rgb_reg = 3'b101; end
            18'b111000011101010100: begin rgb_reg = 3'b101; end
            18'b111000011101010111: begin rgb_reg = 3'b101; end
            18'b111000011101011000: begin rgb_reg = 3'b101; end
            18'b111000011101100000: begin rgb_reg = 3'b101; end
            18'b111000011101100001: begin rgb_reg = 3'b101; end
            18'b111000011101101011: begin rgb_reg = 3'b101; end
            18'b111000011101101100: begin rgb_reg = 3'b101; end
            18'b111000011101110010: begin rgb_reg = 3'b101; end
            18'b111000011101110011: begin rgb_reg = 3'b101; end
            18'b111000011101110111: begin rgb_reg = 3'b101; end
            18'b111000011101111000: begin rgb_reg = 3'b101; end
            18'b111000011101111011: begin rgb_reg = 3'b101; end
            18'b111000011101111100: begin rgb_reg = 3'b101; end
            18'b111000011110000000: begin rgb_reg = 3'b101; end
            18'b111000011110000001: begin rgb_reg = 3'b101; end
            18'b111000011110001001: begin rgb_reg = 3'b101; end
            18'b111000011110001010: begin rgb_reg = 3'b101; end
            18'b111000011110001101: begin rgb_reg = 3'b101; end
            18'b111000011110001110: begin rgb_reg = 3'b101; end
            18'b111000011110001111: begin rgb_reg = 3'b101; end
            18'b111000011110010000: begin rgb_reg = 3'b101; end
            18'b111000011110010001: begin rgb_reg = 3'b101; end
            18'b111000011110010010: begin rgb_reg = 3'b101; end
            18'b111000011110010011: begin rgb_reg = 3'b101; end
            18'b111000100001101001: begin rgb_reg = 3'b101; end
            18'b111000100001101010: begin rgb_reg = 3'b101; end
            18'b111000100001101011: begin rgb_reg = 3'b101; end
            18'b111000100001101100: begin rgb_reg = 3'b101; end
            18'b111000100001101101: begin rgb_reg = 3'b101; end
            18'b111000100001101110: begin rgb_reg = 3'b101; end
            18'b111000100001101111: begin rgb_reg = 3'b101; end
            18'b111000100001110000: begin rgb_reg = 3'b101; end
            18'b111000100001110001: begin rgb_reg = 3'b101; end
            18'b111000100001110010: begin rgb_reg = 3'b101; end
            18'b111000100001110011: begin rgb_reg = 3'b101; end
            18'b111000100001111000: begin rgb_reg = 3'b101; end
            18'b111000100001111001: begin rgb_reg = 3'b101; end
            18'b111000100010000100: begin rgb_reg = 3'b101; end
            18'b111000100010000101: begin rgb_reg = 3'b101; end
            18'b111000100010011010: begin rgb_reg = 3'b101; end
            18'b111000100010011011: begin rgb_reg = 3'b101; end
            18'b111000100010011100: begin rgb_reg = 3'b101; end
            18'b111000100010011101: begin rgb_reg = 3'b101; end
            18'b111000100010011110: begin rgb_reg = 3'b101; end
            18'b111000100010011111: begin rgb_reg = 3'b101; end
            18'b111000100010100101: begin rgb_reg = 3'b101; end
            18'b111000100010100110: begin rgb_reg = 3'b101; end
            18'b111000100010100111: begin rgb_reg = 3'b101; end
            18'b111000100010101000: begin rgb_reg = 3'b101; end
            18'b111000100010101001: begin rgb_reg = 3'b101; end
            18'b111000100010101010: begin rgb_reg = 3'b101; end
            18'b111000100010101011: begin rgb_reg = 3'b101; end
            18'b111000100010101100: begin rgb_reg = 3'b101; end
            18'b111000100010101101: begin rgb_reg = 3'b101; end
            18'b111000100010110011: begin rgb_reg = 3'b101; end
            18'b111000100010110100: begin rgb_reg = 3'b101; end
            18'b111000100010110101: begin rgb_reg = 3'b101; end
            18'b111000100010110110: begin rgb_reg = 3'b101; end
            18'b111000100010110111: begin rgb_reg = 3'b101; end
            18'b111000100010111000: begin rgb_reg = 3'b101; end
            18'b111000100010111001: begin rgb_reg = 3'b101; end
            18'b111000100010111010: begin rgb_reg = 3'b101; end
            18'b111000100010111011: begin rgb_reg = 3'b101; end
            18'b111000100010111100: begin rgb_reg = 3'b101; end
            18'b111000100010111101: begin rgb_reg = 3'b101; end
            18'b111000100011000000: begin rgb_reg = 3'b101; end
            18'b111000100011000001: begin rgb_reg = 3'b101; end
            18'b111000100011001110: begin rgb_reg = 3'b101; end
            18'b111000100011001111: begin rgb_reg = 3'b101; end
            18'b111000100011010000: begin rgb_reg = 3'b101; end
            18'b111000100011010001: begin rgb_reg = 3'b101; end
            18'b111000100011010010: begin rgb_reg = 3'b101; end
            18'b111000100011010011: begin rgb_reg = 3'b101; end
            18'b111000100011100000: begin rgb_reg = 3'b101; end
            18'b111000100011100001: begin rgb_reg = 3'b101; end
            18'b111000100011100010: begin rgb_reg = 3'b101; end
            18'b111000100011100011: begin rgb_reg = 3'b101; end
            18'b111000100011100100: begin rgb_reg = 3'b101; end
            18'b111000100011100101: begin rgb_reg = 3'b101; end
            18'b111000100011100110: begin rgb_reg = 3'b101; end
            18'b111000100011100111: begin rgb_reg = 3'b101; end
            18'b111000100011101101: begin rgb_reg = 3'b101; end
            18'b111000100011101110: begin rgb_reg = 3'b101; end
            18'b111000100011101111: begin rgb_reg = 3'b101; end
            18'b111000100011110000: begin rgb_reg = 3'b101; end
            18'b111000100011110001: begin rgb_reg = 3'b101; end
            18'b111000100011110010: begin rgb_reg = 3'b101; end
            18'b111000100011110011: begin rgb_reg = 3'b101; end
            18'b111000100011110100: begin rgb_reg = 3'b101; end
            18'b111000100011110101: begin rgb_reg = 3'b101; end
            18'b111000100011110110: begin rgb_reg = 3'b101; end
            18'b111000100011110111: begin rgb_reg = 3'b101; end
            18'b111000100011111011: begin rgb_reg = 3'b101; end
            18'b111000100011111100: begin rgb_reg = 3'b101; end
            18'b111000100011111101: begin rgb_reg = 3'b101; end
            18'b111000100011111110: begin rgb_reg = 3'b101; end
            18'b111000100011111111: begin rgb_reg = 3'b101; end
            18'b111000100100000000: begin rgb_reg = 3'b101; end
            18'b111000100100000001: begin rgb_reg = 3'b101; end
            18'b111000100100000010: begin rgb_reg = 3'b101; end
            18'b111000100100011000: begin rgb_reg = 3'b101; end
            18'b111000100100011001: begin rgb_reg = 3'b101; end
            18'b111000100100100001: begin rgb_reg = 3'b101; end
            18'b111000100100100010: begin rgb_reg = 3'b101; end
            18'b111000100100101010: begin rgb_reg = 3'b101; end
            18'b111000100100101011: begin rgb_reg = 3'b101; end
            18'b111000100100110011: begin rgb_reg = 3'b101; end
            18'b111000100100110100: begin rgb_reg = 3'b101; end
            18'b111000100101000001: begin rgb_reg = 3'b101; end
            18'b111000100101000010: begin rgb_reg = 3'b101; end
            18'b111000100101001010: begin rgb_reg = 3'b101; end
            18'b111000100101001011: begin rgb_reg = 3'b101; end
            18'b111000100101001110: begin rgb_reg = 3'b101; end
            18'b111000100101001111: begin rgb_reg = 3'b101; end
            18'b111000100101010011: begin rgb_reg = 3'b101; end
            18'b111000100101010111: begin rgb_reg = 3'b101; end
            18'b111000100101011000: begin rgb_reg = 3'b101; end
            18'b111000100101100000: begin rgb_reg = 3'b101; end
            18'b111000100101100001: begin rgb_reg = 3'b101; end
            18'b111000100101101011: begin rgb_reg = 3'b101; end
            18'b111000100101101100: begin rgb_reg = 3'b101; end
            18'b111000100101110010: begin rgb_reg = 3'b101; end
            18'b111000100101110011: begin rgb_reg = 3'b101; end
            18'b111000100101110111: begin rgb_reg = 3'b101; end
            18'b111000100101111011: begin rgb_reg = 3'b101; end
            18'b111000100101111100: begin rgb_reg = 3'b101; end
            18'b111000100110000000: begin rgb_reg = 3'b101; end
            18'b111000100110000001: begin rgb_reg = 3'b101; end
            18'b111000100110001001: begin rgb_reg = 3'b101; end
            18'b111000100110001010: begin rgb_reg = 3'b101; end
            18'b111000100110001101: begin rgb_reg = 3'b101; end
            18'b111000100110001110: begin rgb_reg = 3'b101; end
            18'b111000100110001111: begin rgb_reg = 3'b101; end
            18'b111000100110010000: begin rgb_reg = 3'b101; end
            18'b111000100110010001: begin rgb_reg = 3'b101; end
            18'b111000100110010010: begin rgb_reg = 3'b101; end
            18'b111000101001101001: begin rgb_reg = 3'b101; end
            18'b111000101001101010: begin rgb_reg = 3'b101; end
            18'b111000101001110010: begin rgb_reg = 3'b101; end
            18'b111000101001110011: begin rgb_reg = 3'b101; end
            18'b111000101001111000: begin rgb_reg = 3'b101; end
            18'b111000101001111001: begin rgb_reg = 3'b101; end
            18'b111000101010000100: begin rgb_reg = 3'b101; end
            18'b111000101010000101: begin rgb_reg = 3'b101; end
            18'b111000101010100001: begin rgb_reg = 3'b101; end
            18'b111000101010100010: begin rgb_reg = 3'b101; end
            18'b111000101010100101: begin rgb_reg = 3'b101; end
            18'b111000101010100110: begin rgb_reg = 3'b101; end
            18'b111000101010110011: begin rgb_reg = 3'b101; end
            18'b111000101010110100: begin rgb_reg = 3'b101; end
            18'b111000101010111100: begin rgb_reg = 3'b101; end
            18'b111000101010111101: begin rgb_reg = 3'b101; end
            18'b111000101011000000: begin rgb_reg = 3'b101; end
            18'b111000101011000001: begin rgb_reg = 3'b101; end
            18'b111000101011001110: begin rgb_reg = 3'b101; end
            18'b111000101011001111: begin rgb_reg = 3'b101; end
            18'b111000101011100000: begin rgb_reg = 3'b101; end
            18'b111000101011100001: begin rgb_reg = 3'b101; end
            18'b111000101011101001: begin rgb_reg = 3'b101; end
            18'b111000101011101010: begin rgb_reg = 3'b101; end
            18'b111000101011101101: begin rgb_reg = 3'b101; end
            18'b111000101011101110: begin rgb_reg = 3'b101; end
            18'b111000101011110110: begin rgb_reg = 3'b101; end
            18'b111000101011110111: begin rgb_reg = 3'b101; end
            18'b111000101011111011: begin rgb_reg = 3'b101; end
            18'b111000101011111100: begin rgb_reg = 3'b101; end
            18'b111000101100000100: begin rgb_reg = 3'b101; end
            18'b111000101100000101: begin rgb_reg = 3'b101; end
            18'b111000101100011000: begin rgb_reg = 3'b101; end
            18'b111000101100011001: begin rgb_reg = 3'b101; end
            18'b111000101100100001: begin rgb_reg = 3'b101; end
            18'b111000101100100010: begin rgb_reg = 3'b101; end
            18'b111000101100101010: begin rgb_reg = 3'b101; end
            18'b111000101100101011: begin rgb_reg = 3'b101; end
            18'b111000101100110011: begin rgb_reg = 3'b101; end
            18'b111000101100110100: begin rgb_reg = 3'b101; end
            18'b111000101101000001: begin rgb_reg = 3'b101; end
            18'b111000101101000010: begin rgb_reg = 3'b101; end
            18'b111000101101001010: begin rgb_reg = 3'b101; end
            18'b111000101101001011: begin rgb_reg = 3'b101; end
            18'b111000101101001110: begin rgb_reg = 3'b101; end
            18'b111000101101001111: begin rgb_reg = 3'b101; end
            18'b111000101101010101: begin rgb_reg = 3'b101; end
            18'b111000101101010110: begin rgb_reg = 3'b101; end
            18'b111000101101010111: begin rgb_reg = 3'b101; end
            18'b111000101101011000: begin rgb_reg = 3'b101; end
            18'b111000101101100000: begin rgb_reg = 3'b101; end
            18'b111000101101100001: begin rgb_reg = 3'b101; end
            18'b111000101101101011: begin rgb_reg = 3'b101; end
            18'b111000101101101100: begin rgb_reg = 3'b101; end
            18'b111000101101110010: begin rgb_reg = 3'b101; end
            18'b111000101101110011: begin rgb_reg = 3'b101; end
            18'b111000101101111001: begin rgb_reg = 3'b101; end
            18'b111000101101111010: begin rgb_reg = 3'b101; end
            18'b111000101101111011: begin rgb_reg = 3'b101; end
            18'b111000101101111100: begin rgb_reg = 3'b101; end
            18'b111000101110000000: begin rgb_reg = 3'b101; end
            18'b111000101110000001: begin rgb_reg = 3'b101; end
            18'b111000101110001001: begin rgb_reg = 3'b101; end
            18'b111000101110001010: begin rgb_reg = 3'b101; end
            18'b111000101110001101: begin rgb_reg = 3'b101; end
            18'b111000101110001110: begin rgb_reg = 3'b101; end
            18'b111000110001101001: begin rgb_reg = 3'b101; end
            18'b111000110001101010: begin rgb_reg = 3'b101; end
            18'b111000110001110010: begin rgb_reg = 3'b101; end
            18'b111000110001110011: begin rgb_reg = 3'b101; end
            18'b111000110001111000: begin rgb_reg = 3'b101; end
            18'b111000110001111001: begin rgb_reg = 3'b101; end
            18'b111000110010000100: begin rgb_reg = 3'b101; end
            18'b111000110010000101: begin rgb_reg = 3'b101; end
            18'b111000110010100001: begin rgb_reg = 3'b101; end
            18'b111000110010100010: begin rgb_reg = 3'b101; end
            18'b111000110010100101: begin rgb_reg = 3'b101; end
            18'b111000110010100110: begin rgb_reg = 3'b101; end
            18'b111000110010110011: begin rgb_reg = 3'b101; end
            18'b111000110010110100: begin rgb_reg = 3'b101; end
            18'b111000110010111100: begin rgb_reg = 3'b101; end
            18'b111000110010111101: begin rgb_reg = 3'b101; end
            18'b111000110011000000: begin rgb_reg = 3'b101; end
            18'b111000110011000001: begin rgb_reg = 3'b101; end
            18'b111000110011001110: begin rgb_reg = 3'b101; end
            18'b111000110011001111: begin rgb_reg = 3'b101; end
            18'b111000110011100000: begin rgb_reg = 3'b101; end
            18'b111000110011100001: begin rgb_reg = 3'b101; end
            18'b111000110011101001: begin rgb_reg = 3'b101; end
            18'b111000110011101010: begin rgb_reg = 3'b101; end
            18'b111000110011101101: begin rgb_reg = 3'b101; end
            18'b111000110011101110: begin rgb_reg = 3'b101; end
            18'b111000110011110110: begin rgb_reg = 3'b101; end
            18'b111000110011110111: begin rgb_reg = 3'b101; end
            18'b111000110011111011: begin rgb_reg = 3'b101; end
            18'b111000110011111100: begin rgb_reg = 3'b101; end
            18'b111000110100000100: begin rgb_reg = 3'b101; end
            18'b111000110100000101: begin rgb_reg = 3'b101; end
            18'b111000110100011000: begin rgb_reg = 3'b101; end
            18'b111000110100011001: begin rgb_reg = 3'b101; end
            18'b111000110100100001: begin rgb_reg = 3'b101; end
            18'b111000110100100010: begin rgb_reg = 3'b101; end
            18'b111000110100101010: begin rgb_reg = 3'b101; end
            18'b111000110100101011: begin rgb_reg = 3'b101; end
            18'b111000110100110011: begin rgb_reg = 3'b101; end
            18'b111000110100110100: begin rgb_reg = 3'b101; end
            18'b111000110101000001: begin rgb_reg = 3'b101; end
            18'b111000110101000010: begin rgb_reg = 3'b101; end
            18'b111000110101001010: begin rgb_reg = 3'b101; end
            18'b111000110101001011: begin rgb_reg = 3'b101; end
            18'b111000110101001110: begin rgb_reg = 3'b101; end
            18'b111000110101001111: begin rgb_reg = 3'b101; end
            18'b111000110101010101: begin rgb_reg = 3'b101; end
            18'b111000110101010110: begin rgb_reg = 3'b101; end
            18'b111000110101010111: begin rgb_reg = 3'b101; end
            18'b111000110101011000: begin rgb_reg = 3'b101; end
            18'b111000110101100000: begin rgb_reg = 3'b101; end
            18'b111000110101100001: begin rgb_reg = 3'b101; end
            18'b111000110101101011: begin rgb_reg = 3'b101; end
            18'b111000110101101100: begin rgb_reg = 3'b101; end
            18'b111000110101110010: begin rgb_reg = 3'b101; end
            18'b111000110101110011: begin rgb_reg = 3'b101; end
            18'b111000110101111001: begin rgb_reg = 3'b101; end
            18'b111000110101111010: begin rgb_reg = 3'b101; end
            18'b111000110101111011: begin rgb_reg = 3'b101; end
            18'b111000110101111100: begin rgb_reg = 3'b101; end
            18'b111000110110000000: begin rgb_reg = 3'b101; end
            18'b111000110110000001: begin rgb_reg = 3'b101; end
            18'b111000110110001001: begin rgb_reg = 3'b101; end
            18'b111000110110001010: begin rgb_reg = 3'b101; end
            18'b111000110110001101: begin rgb_reg = 3'b101; end
            18'b111000110110001110: begin rgb_reg = 3'b101; end
            18'b111000111001101001: begin rgb_reg = 3'b101; end
            18'b111000111001101010: begin rgb_reg = 3'b101; end
            18'b111000111001110010: begin rgb_reg = 3'b101; end
            18'b111000111001110011: begin rgb_reg = 3'b101; end
            18'b111000111001111000: begin rgb_reg = 3'b101; end
            18'b111000111001111001: begin rgb_reg = 3'b101; end
            18'b111000111010000100: begin rgb_reg = 3'b101; end
            18'b111000111010000101: begin rgb_reg = 3'b101; end
            18'b111000111010100001: begin rgb_reg = 3'b101; end
            18'b111000111010100010: begin rgb_reg = 3'b101; end
            18'b111000111010100101: begin rgb_reg = 3'b101; end
            18'b111000111010100110: begin rgb_reg = 3'b101; end
            18'b111000111010110011: begin rgb_reg = 3'b101; end
            18'b111000111010110100: begin rgb_reg = 3'b101; end
            18'b111000111010111100: begin rgb_reg = 3'b101; end
            18'b111000111010111101: begin rgb_reg = 3'b101; end
            18'b111000111011000000: begin rgb_reg = 3'b101; end
            18'b111000111011000001: begin rgb_reg = 3'b101; end
            18'b111000111011001110: begin rgb_reg = 3'b101; end
            18'b111000111011001111: begin rgb_reg = 3'b101; end
            18'b111000111011100000: begin rgb_reg = 3'b101; end
            18'b111000111011100001: begin rgb_reg = 3'b101; end
            18'b111000111011101001: begin rgb_reg = 3'b101; end
            18'b111000111011101010: begin rgb_reg = 3'b101; end
            18'b111000111011101101: begin rgb_reg = 3'b101; end
            18'b111000111011101110: begin rgb_reg = 3'b101; end
            18'b111000111011110110: begin rgb_reg = 3'b101; end
            18'b111000111011110111: begin rgb_reg = 3'b101; end
            18'b111000111011111011: begin rgb_reg = 3'b101; end
            18'b111000111011111100: begin rgb_reg = 3'b101; end
            18'b111000111100000100: begin rgb_reg = 3'b101; end
            18'b111000111100000101: begin rgb_reg = 3'b101; end
            18'b111000111100011000: begin rgb_reg = 3'b101; end
            18'b111000111100011001: begin rgb_reg = 3'b101; end
            18'b111000111100100001: begin rgb_reg = 3'b101; end
            18'b111000111100100010: begin rgb_reg = 3'b101; end
            18'b111000111100101010: begin rgb_reg = 3'b101; end
            18'b111000111100101011: begin rgb_reg = 3'b101; end
            18'b111000111100110011: begin rgb_reg = 3'b101; end
            18'b111000111100110100: begin rgb_reg = 3'b101; end
            18'b111000111101000001: begin rgb_reg = 3'b101; end
            18'b111000111101000010: begin rgb_reg = 3'b101; end
            18'b111000111101001010: begin rgb_reg = 3'b101; end
            18'b111000111101001011: begin rgb_reg = 3'b101; end
            18'b111000111101001110: begin rgb_reg = 3'b101; end
            18'b111000111101001111: begin rgb_reg = 3'b101; end
            18'b111000111101010111: begin rgb_reg = 3'b101; end
            18'b111000111101011000: begin rgb_reg = 3'b101; end
            18'b111000111101100000: begin rgb_reg = 3'b101; end
            18'b111000111101100001: begin rgb_reg = 3'b101; end
            18'b111000111101101011: begin rgb_reg = 3'b101; end
            18'b111000111101101100: begin rgb_reg = 3'b101; end
            18'b111000111101110010: begin rgb_reg = 3'b101; end
            18'b111000111101110011: begin rgb_reg = 3'b101; end
            18'b111000111101111011: begin rgb_reg = 3'b101; end
            18'b111000111101111100: begin rgb_reg = 3'b101; end
            18'b111000111110000000: begin rgb_reg = 3'b101; end
            18'b111000111110000001: begin rgb_reg = 3'b101; end
            18'b111000111110001001: begin rgb_reg = 3'b101; end
            18'b111000111110001010: begin rgb_reg = 3'b101; end
            18'b111000111110001101: begin rgb_reg = 3'b101; end
            18'b111000111110001110: begin rgb_reg = 3'b101; end
            18'b111001000001101001: begin rgb_reg = 3'b101; end
            18'b111001000001101010: begin rgb_reg = 3'b101; end
            18'b111001000001110010: begin rgb_reg = 3'b101; end
            18'b111001000001110011: begin rgb_reg = 3'b101; end
            18'b111001000001111000: begin rgb_reg = 3'b101; end
            18'b111001000001111001: begin rgb_reg = 3'b101; end
            18'b111001000010000100: begin rgb_reg = 3'b101; end
            18'b111001000010000101: begin rgb_reg = 3'b101; end
            18'b111001000010100001: begin rgb_reg = 3'b101; end
            18'b111001000010100010: begin rgb_reg = 3'b101; end
            18'b111001000010100101: begin rgb_reg = 3'b101; end
            18'b111001000010100110: begin rgb_reg = 3'b101; end
            18'b111001000010110011: begin rgb_reg = 3'b101; end
            18'b111001000010110100: begin rgb_reg = 3'b101; end
            18'b111001000010111100: begin rgb_reg = 3'b101; end
            18'b111001000010111101: begin rgb_reg = 3'b101; end
            18'b111001000011000000: begin rgb_reg = 3'b101; end
            18'b111001000011000001: begin rgb_reg = 3'b101; end
            18'b111001000011001110: begin rgb_reg = 3'b101; end
            18'b111001000011001111: begin rgb_reg = 3'b101; end
            18'b111001000011100000: begin rgb_reg = 3'b101; end
            18'b111001000011100001: begin rgb_reg = 3'b101; end
            18'b111001000011101001: begin rgb_reg = 3'b101; end
            18'b111001000011101010: begin rgb_reg = 3'b101; end
            18'b111001000011101101: begin rgb_reg = 3'b101; end
            18'b111001000011101110: begin rgb_reg = 3'b101; end
            18'b111001000011110110: begin rgb_reg = 3'b101; end
            18'b111001000011110111: begin rgb_reg = 3'b101; end
            18'b111001000011111011: begin rgb_reg = 3'b101; end
            18'b111001000011111100: begin rgb_reg = 3'b101; end
            18'b111001000100000100: begin rgb_reg = 3'b101; end
            18'b111001000100000101: begin rgb_reg = 3'b101; end
            18'b111001000100011000: begin rgb_reg = 3'b101; end
            18'b111001000100011001: begin rgb_reg = 3'b101; end
            18'b111001000100100001: begin rgb_reg = 3'b101; end
            18'b111001000100100010: begin rgb_reg = 3'b101; end
            18'b111001000100101010: begin rgb_reg = 3'b101; end
            18'b111001000100101011: begin rgb_reg = 3'b101; end
            18'b111001000100110011: begin rgb_reg = 3'b101; end
            18'b111001000100110100: begin rgb_reg = 3'b101; end
            18'b111001000101000001: begin rgb_reg = 3'b101; end
            18'b111001000101000010: begin rgb_reg = 3'b101; end
            18'b111001000101001010: begin rgb_reg = 3'b101; end
            18'b111001000101001011: begin rgb_reg = 3'b101; end
            18'b111001000101001110: begin rgb_reg = 3'b101; end
            18'b111001000101001111: begin rgb_reg = 3'b101; end
            18'b111001000101010111: begin rgb_reg = 3'b101; end
            18'b111001000101011000: begin rgb_reg = 3'b101; end
            18'b111001000101100000: begin rgb_reg = 3'b101; end
            18'b111001000101100001: begin rgb_reg = 3'b101; end
            18'b111001000101101011: begin rgb_reg = 3'b101; end
            18'b111001000101101100: begin rgb_reg = 3'b101; end
            18'b111001000101110010: begin rgb_reg = 3'b101; end
            18'b111001000101110011: begin rgb_reg = 3'b101; end
            18'b111001000101111011: begin rgb_reg = 3'b101; end
            18'b111001000101111100: begin rgb_reg = 3'b101; end
            18'b111001000110000000: begin rgb_reg = 3'b101; end
            18'b111001000110000001: begin rgb_reg = 3'b101; end
            18'b111001000110001001: begin rgb_reg = 3'b101; end
            18'b111001000110001010: begin rgb_reg = 3'b101; end
            18'b111001000110001101: begin rgb_reg = 3'b101; end
            18'b111001000110001110: begin rgb_reg = 3'b101; end
            18'b111001001001101001: begin rgb_reg = 3'b101; end
            18'b111001001001101010: begin rgb_reg = 3'b101; end
            18'b111001001001110010: begin rgb_reg = 3'b101; end
            18'b111001001001110011: begin rgb_reg = 3'b101; end
            18'b111001001001111000: begin rgb_reg = 3'b101; end
            18'b111001001001111001: begin rgb_reg = 3'b101; end
            18'b111001001010000100: begin rgb_reg = 3'b101; end
            18'b111001001010000101: begin rgb_reg = 3'b101; end
            18'b111001001010011000: begin rgb_reg = 3'b101; end
            18'b111001001010011001: begin rgb_reg = 3'b101; end
            18'b111001001010100001: begin rgb_reg = 3'b101; end
            18'b111001001010100010: begin rgb_reg = 3'b101; end
            18'b111001001010100101: begin rgb_reg = 3'b101; end
            18'b111001001010100110: begin rgb_reg = 3'b101; end
            18'b111001001010110011: begin rgb_reg = 3'b101; end
            18'b111001001010110100: begin rgb_reg = 3'b101; end
            18'b111001001010111100: begin rgb_reg = 3'b101; end
            18'b111001001010111101: begin rgb_reg = 3'b101; end
            18'b111001001011000000: begin rgb_reg = 3'b101; end
            18'b111001001011000001: begin rgb_reg = 3'b101; end
            18'b111001001011001010: begin rgb_reg = 3'b101; end
            18'b111001001011001110: begin rgb_reg = 3'b101; end
            18'b111001001011001111: begin rgb_reg = 3'b101; end
            18'b111001001011100000: begin rgb_reg = 3'b101; end
            18'b111001001011100001: begin rgb_reg = 3'b101; end
            18'b111001001011101001: begin rgb_reg = 3'b101; end
            18'b111001001011101010: begin rgb_reg = 3'b101; end
            18'b111001001011101101: begin rgb_reg = 3'b101; end
            18'b111001001011101110: begin rgb_reg = 3'b101; end
            18'b111001001011110110: begin rgb_reg = 3'b101; end
            18'b111001001011110111: begin rgb_reg = 3'b101; end
            18'b111001001011111011: begin rgb_reg = 3'b101; end
            18'b111001001011111100: begin rgb_reg = 3'b101; end
            18'b111001001100000100: begin rgb_reg = 3'b101; end
            18'b111001001100000101: begin rgb_reg = 3'b101; end
            18'b111001001100011000: begin rgb_reg = 3'b101; end
            18'b111001001100011001: begin rgb_reg = 3'b101; end
            18'b111001001100100001: begin rgb_reg = 3'b101; end
            18'b111001001100100010: begin rgb_reg = 3'b101; end
            18'b111001001100101010: begin rgb_reg = 3'b101; end
            18'b111001001100101011: begin rgb_reg = 3'b101; end
            18'b111001001100110011: begin rgb_reg = 3'b101; end
            18'b111001001100110100: begin rgb_reg = 3'b101; end
            18'b111001001100111100: begin rgb_reg = 3'b101; end
            18'b111001001100111101: begin rgb_reg = 3'b101; end
            18'b111001001101000001: begin rgb_reg = 3'b101; end
            18'b111001001101000010: begin rgb_reg = 3'b101; end
            18'b111001001101001010: begin rgb_reg = 3'b101; end
            18'b111001001101001011: begin rgb_reg = 3'b101; end
            18'b111001001101001110: begin rgb_reg = 3'b101; end
            18'b111001001101001111: begin rgb_reg = 3'b101; end
            18'b111001001101010111: begin rgb_reg = 3'b101; end
            18'b111001001101011000: begin rgb_reg = 3'b101; end
            18'b111001001101100000: begin rgb_reg = 3'b101; end
            18'b111001001101100001: begin rgb_reg = 3'b101; end
            18'b111001001101101011: begin rgb_reg = 3'b101; end
            18'b111001001101101100: begin rgb_reg = 3'b101; end
            18'b111001001101110010: begin rgb_reg = 3'b101; end
            18'b111001001101110011: begin rgb_reg = 3'b101; end
            18'b111001001101111011: begin rgb_reg = 3'b101; end
            18'b111001001101111100: begin rgb_reg = 3'b101; end
            18'b111001001110000000: begin rgb_reg = 3'b101; end
            18'b111001001110000001: begin rgb_reg = 3'b101; end
            18'b111001001110001001: begin rgb_reg = 3'b101; end
            18'b111001001110001010: begin rgb_reg = 3'b101; end
            18'b111001001110001101: begin rgb_reg = 3'b101; end
            18'b111001001110001110: begin rgb_reg = 3'b101; end
            18'b111001010001101001: begin rgb_reg = 3'b101; end
            18'b111001010001101010: begin rgb_reg = 3'b101; end
            18'b111001010001110010: begin rgb_reg = 3'b101; end
            18'b111001010001110011: begin rgb_reg = 3'b101; end
            18'b111001010001111000: begin rgb_reg = 3'b101; end
            18'b111001010001111001: begin rgb_reg = 3'b101; end
            18'b111001010010000100: begin rgb_reg = 3'b101; end
            18'b111001010010000101: begin rgb_reg = 3'b101; end
            18'b111001010010011000: begin rgb_reg = 3'b101; end
            18'b111001010010011001: begin rgb_reg = 3'b101; end
            18'b111001010010100001: begin rgb_reg = 3'b101; end
            18'b111001010010100010: begin rgb_reg = 3'b101; end
            18'b111001010010100101: begin rgb_reg = 3'b101; end
            18'b111001010010100110: begin rgb_reg = 3'b101; end
            18'b111001010010110011: begin rgb_reg = 3'b101; end
            18'b111001010010110100: begin rgb_reg = 3'b101; end
            18'b111001010010111100: begin rgb_reg = 3'b101; end
            18'b111001010010111101: begin rgb_reg = 3'b101; end
            18'b111001010011000000: begin rgb_reg = 3'b101; end
            18'b111001010011000001: begin rgb_reg = 3'b101; end
            18'b111001010011001001: begin rgb_reg = 3'b101; end
            18'b111001010011001010: begin rgb_reg = 3'b101; end
            18'b111001010011001110: begin rgb_reg = 3'b101; end
            18'b111001010011001111: begin rgb_reg = 3'b101; end
            18'b111001010011100000: begin rgb_reg = 3'b101; end
            18'b111001010011100001: begin rgb_reg = 3'b101; end
            18'b111001010011101001: begin rgb_reg = 3'b101; end
            18'b111001010011101010: begin rgb_reg = 3'b101; end
            18'b111001010011101101: begin rgb_reg = 3'b101; end
            18'b111001010011101110: begin rgb_reg = 3'b101; end
            18'b111001010011110110: begin rgb_reg = 3'b101; end
            18'b111001010011110111: begin rgb_reg = 3'b101; end
            18'b111001010011111011: begin rgb_reg = 3'b101; end
            18'b111001010011111100: begin rgb_reg = 3'b101; end
            18'b111001010100000100: begin rgb_reg = 3'b101; end
            18'b111001010100000101: begin rgb_reg = 3'b101; end
            18'b111001010100011000: begin rgb_reg = 3'b101; end
            18'b111001010100011001: begin rgb_reg = 3'b101; end
            18'b111001010100100001: begin rgb_reg = 3'b101; end
            18'b111001010100100010: begin rgb_reg = 3'b101; end
            18'b111001010100101010: begin rgb_reg = 3'b101; end
            18'b111001010100101011: begin rgb_reg = 3'b101; end
            18'b111001010100110011: begin rgb_reg = 3'b101; end
            18'b111001010100110100: begin rgb_reg = 3'b101; end
            18'b111001010100111100: begin rgb_reg = 3'b101; end
            18'b111001010100111101: begin rgb_reg = 3'b101; end
            18'b111001010101000001: begin rgb_reg = 3'b101; end
            18'b111001010101000010: begin rgb_reg = 3'b101; end
            18'b111001010101001010: begin rgb_reg = 3'b101; end
            18'b111001010101001011: begin rgb_reg = 3'b101; end
            18'b111001010101001110: begin rgb_reg = 3'b101; end
            18'b111001010101001111: begin rgb_reg = 3'b101; end
            18'b111001010101010111: begin rgb_reg = 3'b101; end
            18'b111001010101011000: begin rgb_reg = 3'b101; end
            18'b111001010101100000: begin rgb_reg = 3'b101; end
            18'b111001010101100001: begin rgb_reg = 3'b101; end
            18'b111001010101101011: begin rgb_reg = 3'b101; end
            18'b111001010101101100: begin rgb_reg = 3'b101; end
            18'b111001010101110010: begin rgb_reg = 3'b101; end
            18'b111001010101110011: begin rgb_reg = 3'b101; end
            18'b111001010101111011: begin rgb_reg = 3'b101; end
            18'b111001010101111100: begin rgb_reg = 3'b101; end
            18'b111001010110000000: begin rgb_reg = 3'b101; end
            18'b111001010110000001: begin rgb_reg = 3'b101; end
            18'b111001010110001001: begin rgb_reg = 3'b101; end
            18'b111001010110001010: begin rgb_reg = 3'b101; end
            18'b111001010110001101: begin rgb_reg = 3'b101; end
            18'b111001010110001110: begin rgb_reg = 3'b101; end
            18'b111001011001101001: begin rgb_reg = 3'b101; end
            18'b111001011001101010: begin rgb_reg = 3'b101; end
            18'b111001011001110010: begin rgb_reg = 3'b101; end
            18'b111001011001110011: begin rgb_reg = 3'b101; end
            18'b111001011001111000: begin rgb_reg = 3'b101; end
            18'b111001011001111001: begin rgb_reg = 3'b101; end
            18'b111001011001111010: begin rgb_reg = 3'b101; end
            18'b111001011010000100: begin rgb_reg = 3'b101; end
            18'b111001011010000101: begin rgb_reg = 3'b101; end
            18'b111001011010100101: begin rgb_reg = 3'b101; end
            18'b111001011010100110: begin rgb_reg = 3'b101; end
            18'b111001011010110011: begin rgb_reg = 3'b101; end
            18'b111001011010110100: begin rgb_reg = 3'b101; end
            18'b111001011010111100: begin rgb_reg = 3'b101; end
            18'b111001011010111101: begin rgb_reg = 3'b101; end
            18'b111001011011001110: begin rgb_reg = 3'b101; end
            18'b111001011011001111: begin rgb_reg = 3'b101; end
            18'b111001011011100000: begin rgb_reg = 3'b101; end
            18'b111001011011100001: begin rgb_reg = 3'b101; end
            18'b111001011011101101: begin rgb_reg = 3'b101; end
            18'b111001011011101110: begin rgb_reg = 3'b101; end
            18'b111001011011110110: begin rgb_reg = 3'b101; end
            18'b111001011011110111: begin rgb_reg = 3'b101; end
            18'b111001011011111011: begin rgb_reg = 3'b101; end
            18'b111001011011111100: begin rgb_reg = 3'b101; end
            18'b111001011100000100: begin rgb_reg = 3'b101; end
            18'b111001011100000101: begin rgb_reg = 3'b101; end
            18'b111001011100011000: begin rgb_reg = 3'b101; end
            18'b111001011100011001: begin rgb_reg = 3'b101; end
            18'b111001011101001110: begin rgb_reg = 3'b101; end
            18'b111001011101001111: begin rgb_reg = 3'b101; end
            18'b111001011101010111: begin rgb_reg = 3'b101; end
            18'b111001011101011000: begin rgb_reg = 3'b101; end
            18'b111001011101100000: begin rgb_reg = 3'b101; end
            18'b111001011101100001: begin rgb_reg = 3'b101; end
            18'b111001011101101011: begin rgb_reg = 3'b101; end
            18'b111001011101101100: begin rgb_reg = 3'b101; end
            18'b111001011101101101: begin rgb_reg = 3'b101; end
            18'b111001011101110010: begin rgb_reg = 3'b101; end
            18'b111001011101110011: begin rgb_reg = 3'b101; end
            18'b111001011101111011: begin rgb_reg = 3'b101; end
            18'b111001011101111100: begin rgb_reg = 3'b101; end
            18'b111001011110001101: begin rgb_reg = 3'b101; end
            18'b111001011110001110: begin rgb_reg = 3'b101; end
            18'b111001100001101001: begin rgb_reg = 3'b101; end
            18'b111001100001101010: begin rgb_reg = 3'b101; end
            18'b111001100001110010: begin rgb_reg = 3'b101; end
            18'b111001100001110011: begin rgb_reg = 3'b101; end
            18'b111001100001110110: begin rgb_reg = 3'b101; end
            18'b111001100001110111: begin rgb_reg = 3'b101; end
            18'b111001100001111000: begin rgb_reg = 3'b101; end
            18'b111001100001111001: begin rgb_reg = 3'b101; end
            18'b111001100001111010: begin rgb_reg = 3'b101; end
            18'b111001100001111011: begin rgb_reg = 3'b101; end
            18'b111001100001111100: begin rgb_reg = 3'b101; end
            18'b111001100010000100: begin rgb_reg = 3'b101; end
            18'b111001100010000101: begin rgb_reg = 3'b101; end
            18'b111001100010011010: begin rgb_reg = 3'b101; end
            18'b111001100010011011: begin rgb_reg = 3'b101; end
            18'b111001100010011100: begin rgb_reg = 3'b101; end
            18'b111001100010011101: begin rgb_reg = 3'b101; end
            18'b111001100010011110: begin rgb_reg = 3'b101; end
            18'b111001100010011111: begin rgb_reg = 3'b101; end
            18'b111001100010100000: begin rgb_reg = 3'b101; end
            18'b111001100010100101: begin rgb_reg = 3'b101; end
            18'b111001100010100110: begin rgb_reg = 3'b101; end
            18'b111001100010110011: begin rgb_reg = 3'b101; end
            18'b111001100010110100: begin rgb_reg = 3'b101; end
            18'b111001100010111100: begin rgb_reg = 3'b101; end
            18'b111001100010111101: begin rgb_reg = 3'b101; end
            18'b111001100011000011: begin rgb_reg = 3'b101; end
            18'b111001100011000100: begin rgb_reg = 3'b101; end
            18'b111001100011000101: begin rgb_reg = 3'b101; end
            18'b111001100011000110: begin rgb_reg = 3'b101; end
            18'b111001100011000111: begin rgb_reg = 3'b101; end
            18'b111001100011001000: begin rgb_reg = 3'b101; end
            18'b111001100011001110: begin rgb_reg = 3'b101; end
            18'b111001100011001111: begin rgb_reg = 3'b101; end
            18'b111001100011010000: begin rgb_reg = 3'b101; end
            18'b111001100011010001: begin rgb_reg = 3'b101; end
            18'b111001100011010010: begin rgb_reg = 3'b101; end
            18'b111001100011010011: begin rgb_reg = 3'b101; end
            18'b111001100011010100: begin rgb_reg = 3'b101; end
            18'b111001100011010101: begin rgb_reg = 3'b101; end
            18'b111001100011010110: begin rgb_reg = 3'b101; end
            18'b111001100011010111: begin rgb_reg = 3'b101; end
            18'b111001100011011000: begin rgb_reg = 3'b101; end
            18'b111001100011100000: begin rgb_reg = 3'b101; end
            18'b111001100011100001: begin rgb_reg = 3'b101; end
            18'b111001100011100010: begin rgb_reg = 3'b101; end
            18'b111001100011100011: begin rgb_reg = 3'b101; end
            18'b111001100011100100: begin rgb_reg = 3'b101; end
            18'b111001100011100101: begin rgb_reg = 3'b101; end
            18'b111001100011100110: begin rgb_reg = 3'b101; end
            18'b111001100011100111: begin rgb_reg = 3'b101; end
            18'b111001100011101000: begin rgb_reg = 3'b101; end
            18'b111001100011101101: begin rgb_reg = 3'b101; end
            18'b111001100011101110: begin rgb_reg = 3'b101; end
            18'b111001100011110110: begin rgb_reg = 3'b101; end
            18'b111001100011110111: begin rgb_reg = 3'b101; end
            18'b111001100011111011: begin rgb_reg = 3'b101; end
            18'b111001100011111100: begin rgb_reg = 3'b101; end
            18'b111001100100000100: begin rgb_reg = 3'b101; end
            18'b111001100100000101: begin rgb_reg = 3'b101; end
            18'b111001100100011000: begin rgb_reg = 3'b101; end
            18'b111001100100011001: begin rgb_reg = 3'b101; end
            18'b111001100100100011: begin rgb_reg = 3'b101; end
            18'b111001100100100100: begin rgb_reg = 3'b101; end
            18'b111001100100100101: begin rgb_reg = 3'b101; end
            18'b111001100100100110: begin rgb_reg = 3'b101; end
            18'b111001100100100111: begin rgb_reg = 3'b101; end
            18'b111001100100101000: begin rgb_reg = 3'b101; end
            18'b111001100100101001: begin rgb_reg = 3'b101; end
            18'b111001100100110101: begin rgb_reg = 3'b101; end
            18'b111001100100110110: begin rgb_reg = 3'b101; end
            18'b111001100100110111: begin rgb_reg = 3'b101; end
            18'b111001100100111000: begin rgb_reg = 3'b101; end
            18'b111001100100111001: begin rgb_reg = 3'b101; end
            18'b111001100100111010: begin rgb_reg = 3'b101; end
            18'b111001100100111011: begin rgb_reg = 3'b101; end
            18'b111001100101000011: begin rgb_reg = 3'b101; end
            18'b111001100101000100: begin rgb_reg = 3'b101; end
            18'b111001100101000101: begin rgb_reg = 3'b101; end
            18'b111001100101000110: begin rgb_reg = 3'b101; end
            18'b111001100101000111: begin rgb_reg = 3'b101; end
            18'b111001100101001000: begin rgb_reg = 3'b101; end
            18'b111001100101001110: begin rgb_reg = 3'b101; end
            18'b111001100101001111: begin rgb_reg = 3'b101; end
            18'b111001100101010111: begin rgb_reg = 3'b101; end
            18'b111001100101011000: begin rgb_reg = 3'b101; end
            18'b111001100101100000: begin rgb_reg = 3'b101; end
            18'b111001100101100001: begin rgb_reg = 3'b101; end
            18'b111001100101101001: begin rgb_reg = 3'b101; end
            18'b111001100101101010: begin rgb_reg = 3'b101; end
            18'b111001100101101011: begin rgb_reg = 3'b101; end
            18'b111001100101101100: begin rgb_reg = 3'b101; end
            18'b111001100101101101: begin rgb_reg = 3'b101; end
            18'b111001100101101110: begin rgb_reg = 3'b101; end
            18'b111001100101101111: begin rgb_reg = 3'b101; end
            18'b111001100101110010: begin rgb_reg = 3'b101; end
            18'b111001100101110011: begin rgb_reg = 3'b101; end
            18'b111001100101111011: begin rgb_reg = 3'b101; end
            18'b111001100101111100: begin rgb_reg = 3'b101; end
            18'b111001100110000010: begin rgb_reg = 3'b101; end
            18'b111001100110000011: begin rgb_reg = 3'b101; end
            18'b111001100110000100: begin rgb_reg = 3'b101; end
            18'b111001100110000101: begin rgb_reg = 3'b101; end
            18'b111001100110000110: begin rgb_reg = 3'b101; end
            18'b111001100110000111: begin rgb_reg = 3'b101; end
            18'b111001100110001101: begin rgb_reg = 3'b101; end
            18'b111001100110001110: begin rgb_reg = 3'b101; end
            18'b111001100110001111: begin rgb_reg = 3'b101; end
            18'b111001100110010000: begin rgb_reg = 3'b101; end
            18'b111001100110010001: begin rgb_reg = 3'b101; end
            18'b111001100110010010: begin rgb_reg = 3'b101; end
            18'b111001100110010011: begin rgb_reg = 3'b101; end
            18'b111001100110010100: begin rgb_reg = 3'b101; end
            18'b111001100110010101: begin rgb_reg = 3'b101; end
            18'b111001100110010110: begin rgb_reg = 3'b101; end
            18'b111001100110010111: begin rgb_reg = 3'b101; end
            18'b111001101001101001: begin rgb_reg = 3'b101; end
            18'b111001101001110010: begin rgb_reg = 3'b101; end
            18'b111001101001110110: begin rgb_reg = 3'b101; end
            18'b111001101001110111: begin rgb_reg = 3'b101; end
            18'b111001101001111000: begin rgb_reg = 3'b101; end
            18'b111001101001111001: begin rgb_reg = 3'b101; end
            18'b111001101001111010: begin rgb_reg = 3'b101; end
            18'b111001101001111011: begin rgb_reg = 3'b101; end
            18'b111001101010000100: begin rgb_reg = 3'b101; end
            18'b111001101010011010: begin rgb_reg = 3'b101; end
            18'b111001101010011011: begin rgb_reg = 3'b101; end
            18'b111001101010011100: begin rgb_reg = 3'b101; end
            18'b111001101010011101: begin rgb_reg = 3'b101; end
            18'b111001101010011110: begin rgb_reg = 3'b101; end
            18'b111001101010011111: begin rgb_reg = 3'b101; end
            18'b111001101010100110: begin rgb_reg = 3'b101; end
            18'b111001101010110011: begin rgb_reg = 3'b101; end
            18'b111001101010110100: begin rgb_reg = 3'b101; end
            18'b111001101010111100: begin rgb_reg = 3'b101; end
            18'b111001101010111101: begin rgb_reg = 3'b101; end
            18'b111001101011000011: begin rgb_reg = 3'b101; end
            18'b111001101011000100: begin rgb_reg = 3'b101; end
            18'b111001101011000101: begin rgb_reg = 3'b101; end
            18'b111001101011000110: begin rgb_reg = 3'b101; end
            18'b111001101011000111: begin rgb_reg = 3'b101; end
            18'b111001101011001000: begin rgb_reg = 3'b101; end
            18'b111001101011001110: begin rgb_reg = 3'b101; end
            18'b111001101011001111: begin rgb_reg = 3'b101; end
            18'b111001101011010000: begin rgb_reg = 3'b101; end
            18'b111001101011010001: begin rgb_reg = 3'b101; end
            18'b111001101011010010: begin rgb_reg = 3'b101; end
            18'b111001101011010011: begin rgb_reg = 3'b101; end
            18'b111001101011010100: begin rgb_reg = 3'b101; end
            18'b111001101011010101: begin rgb_reg = 3'b101; end
            18'b111001101011010110: begin rgb_reg = 3'b101; end
            18'b111001101011010111: begin rgb_reg = 3'b101; end
            18'b111001101011011000: begin rgb_reg = 3'b101; end
            18'b111001101011100000: begin rgb_reg = 3'b101; end
            18'b111001101011100001: begin rgb_reg = 3'b101; end
            18'b111001101011100010: begin rgb_reg = 3'b101; end
            18'b111001101011100011: begin rgb_reg = 3'b101; end
            18'b111001101011100100: begin rgb_reg = 3'b101; end
            18'b111001101011100101: begin rgb_reg = 3'b101; end
            18'b111001101011100110: begin rgb_reg = 3'b101; end
            18'b111001101011100111: begin rgb_reg = 3'b101; end
            18'b111001101011101110: begin rgb_reg = 3'b101; end
            18'b111001101011110111: begin rgb_reg = 3'b101; end
            18'b111001101011111011: begin rgb_reg = 3'b101; end
            18'b111001101011111100: begin rgb_reg = 3'b101; end
            18'b111001101100000100: begin rgb_reg = 3'b101; end
            18'b111001101100000101: begin rgb_reg = 3'b101; end
            18'b111001101100011000: begin rgb_reg = 3'b101; end
            18'b111001101100011001: begin rgb_reg = 3'b101; end
            18'b111001101100100100: begin rgb_reg = 3'b101; end
            18'b111001101100100101: begin rgb_reg = 3'b101; end
            18'b111001101100100110: begin rgb_reg = 3'b101; end
            18'b111001101100100111: begin rgb_reg = 3'b101; end
            18'b111001101100101000: begin rgb_reg = 3'b101; end
            18'b111001101100101001: begin rgb_reg = 3'b101; end
            18'b111001101100110110: begin rgb_reg = 3'b101; end
            18'b111001101100110111: begin rgb_reg = 3'b101; end
            18'b111001101100111000: begin rgb_reg = 3'b101; end
            18'b111001101100111001: begin rgb_reg = 3'b101; end
            18'b111001101100111010: begin rgb_reg = 3'b101; end
            18'b111001101100111011: begin rgb_reg = 3'b101; end
            18'b111001101101000011: begin rgb_reg = 3'b101; end
            18'b111001101101000100: begin rgb_reg = 3'b101; end
            18'b111001101101000101: begin rgb_reg = 3'b101; end
            18'b111001101101000110: begin rgb_reg = 3'b101; end
            18'b111001101101000111: begin rgb_reg = 3'b101; end
            18'b111001101101001000: begin rgb_reg = 3'b101; end
            18'b111001101101001110: begin rgb_reg = 3'b101; end
            18'b111001101101001111: begin rgb_reg = 3'b101; end
            18'b111001101101010111: begin rgb_reg = 3'b101; end
            18'b111001101101011000: begin rgb_reg = 3'b101; end
            18'b111001101101100000: begin rgb_reg = 3'b101; end
            18'b111001101101100001: begin rgb_reg = 3'b101; end
            18'b111001101101101001: begin rgb_reg = 3'b101; end
            18'b111001101101101010: begin rgb_reg = 3'b101; end
            18'b111001101101101011: begin rgb_reg = 3'b101; end
            18'b111001101101101100: begin rgb_reg = 3'b101; end
            18'b111001101101101101: begin rgb_reg = 3'b101; end
            18'b111001101101101110: begin rgb_reg = 3'b101; end
            18'b111001101101110010: begin rgb_reg = 3'b101; end
            18'b111001101101110011: begin rgb_reg = 3'b101; end
            18'b111001101101111011: begin rgb_reg = 3'b101; end
            18'b111001101101111100: begin rgb_reg = 3'b101; end
            18'b111001101110000010: begin rgb_reg = 3'b101; end
            18'b111001101110000011: begin rgb_reg = 3'b101; end
            18'b111001101110000100: begin rgb_reg = 3'b101; end
            18'b111001101110000101: begin rgb_reg = 3'b101; end
            18'b111001101110000110: begin rgb_reg = 3'b101; end
            18'b111001101110000111: begin rgb_reg = 3'b101; end
            18'b111001101110001101: begin rgb_reg = 3'b101; end
            18'b111001101110001110: begin rgb_reg = 3'b101; end
            18'b111001101110001111: begin rgb_reg = 3'b101; end
            18'b111001101110010000: begin rgb_reg = 3'b101; end
            18'b111001101110010001: begin rgb_reg = 3'b101; end
            18'b111001101110010010: begin rgb_reg = 3'b101; end
            18'b111001101110010011: begin rgb_reg = 3'b101; end
            18'b111001101110010100: begin rgb_reg = 3'b101; end
            18'b111001101110010101: begin rgb_reg = 3'b101; end
            18'b111001101110010110: begin rgb_reg = 3'b101; end
            18'b111001101110010111: begin rgb_reg = 3'b101; end
            default: begin rgb_reg = 3'b000; end
        endcase
    end  
endmodule
